XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����m���6�� ���{��%�X�C�!��<��������uɏrOh M���b�Jb|M��Gvj���
���	M����j�u���1ϑ(���Xj��S�п�k���ą�Bzq��v5�f"�"i�PP���q�����Ҥn2��vL>(b��p���q8�X�y�t�J#S
X݂:5s���`7���X�����w�+ǅS�&�-��=�/8����Y��S�^z#I
t7~���^���=�s�0{sfd�=^!���)����ʦ��$�
ӣX �%�i�s"@������<�;�7O槔~6�8�m�9h��1G���:D�fq�q2�$KMYf��V��K��KV	�ؔ�
oR_�Tp�o���#-S�l�S��tʘ��3�_}z�ʐ`�V�
����Oה�Y����
���-��5���Y�-��{ڦ�1��c�5�������h�HR��jd6�j�!_da\��{Vb��"�;�����_*`C/;n��o�߷��������G��XU,��ӻ�΅�-��&W��6�1?�>�4�/��1�M���u�R&ނ�"���h�q�1�D�.�&Qy�h�(�8ذ07ET��֥뾪.����0pΈPnB���6�"��f�ea��/�Ʀר���P[�?�`��tR�bqr�?D�}�f#�O6W���*"���ZOK-Ԙ�<��,V)�2ڠϏ%�49���h��ݯd�\iK�97i�Rr�I�DU�y����?����С�XlxVHYEB    6315    1790�l��ӑ:��6�����ohU�u�8a�V`��^�!��>�]$D�Z�p=ړ��8�_�K��R�}��`����춷������ň�ǈK�����(��{� !��<��	�%��Q�S�r��_ZV)���r^~����
�@i�Eձ�x.�-�pꐢ'K)N����6��p�ZpS��,��
�#]Y��ߛJ���WmZ�Z�V�Q�O�i�K��	i�G�n�(�* ZȀ :�=��j����;`��H���x~��m�@5Xn?�QKא��sAD��b`=[���h���?�CP�� ]������L;֓F�X
����&>rᕞ\巚���?j;��{�tx	qW��LJ��Mq��;i�[��%8�"���9���fg�p���k�t�P"K#0���ގ����(��LyM�Jxew{#L�I��^���!��V^�ay�D�N^�A�0")����"��s��1�W�G>�p�82U�6�9 �9-��fm��PV^���(*&"�3��<ڶ������t[*T�
N�q6�Z͂ar��5?�������[8��V:�A�ȫI=��˥����^C��0���Z"	��� ��>�l�r�}J�hq(�S��񲣦Q��@�|s��*S���o$=[=��D"LQ��x��s�n�p�h��i��� ��X�g�E,M���l<��C"�#�vzn&�4�`�������GI�v/�2��R�x\�+��B��^h9�y Y\`f�^��5��=���W1u��\�%r��n�����M\��O�9�Z4:�qzz���F揗
/f�4�Y)�0�=\����䪾M�OJt�BJ�G�� � ��H$U,(���l4�����=����-K-�19B�)�mp���l`�0-PoV����⧿kbM^L����T�MF���{�)�a��k����ٟՠ�ծ��g�5�F0ѣ��s����Y ���}�ޫ��)���b݂��R=�Tڒ޴ %�ti=O�7|�Gr���2-Ԧ�ۤz�U.5�,V9��=��b�/ �����UE:֠sj��*3&%-�-�q�0g��Qh��Pa޴�� ���s}�ù���?���q�V���5�L2�c�"�R��i�⪊>-�G�B۴�� !��C��+n���o��G�\��T'"8��+��.٭��K]�@^bW2㈞(r�vE�	����f�����������^*%;GGp�)�U-�bϙ�}l)iC�Me�IX���@%�(D5�'&��Y�!��߿��5��G��IO��?�������{�iOi�Am��b9���?e��6\u]�;��\כ�D�R���0:�5H�&C���!i�8�HGD�#�і����Xw[�A��jvԭ�� �#p�3}��;�4�j��G䧉
�2�z�Ȝ���8�#q�okX����D����bdD��H�z��b��Fo����z�D��-�$���+�T��U�˾�_TH���6i+�F$��l���)��l1����3S�w�#U>���f�N~�¾����!7vvy�t)��6W��7u��!_�C��]OKˣlU�}�w���E�C'M�X�td���:����]r����n u�tvn5�:�M��0���Nʉر���g�{�#�	 �����ԙ���<H|<�<2?L�} �h�+@	�O�d���B�k���Ct�U�n��#t���D]4~��0a����4l+G��='yKh����4�'t�U��G��M2��c��;zp_�bO��_{~`!#E%L�|��q�z���=�{��&|�����͜��+�h�ژ��hCR z,���\�����Oe
L��1���P����d�;:O�Ԝ�=����
5��j��dٴ�Q[�Mdwn�ީY�ț�	 ��ͳ����|��t��:@�v��߼i�u�Y�t��S�!�Ӫ���,��o��vbd�v��E�0Bj���gP�*b+$eF<�ԍ��rJY"Iζ�=ǳb]�ќX���������ڌZW��2���w5-��-� |�Y2:/+��nD����#EZOU�m�Ё�����)��o��g�>��^�3���p����|�~<l(d��`K���ϸ��K$��+b������r!_��<3�^pB������/Ht�]�ůK��Bʃ��ǜ V�fn=��hj������r��%4�4f���=�a�K���)usZ��n�I�j�V=DQ�=�2n�� �z�s�����K����{o�Y� a(8���Շ6ay�%����?.�~7H�i���_��b{�U��n
�{��ʠ��BD�0���4 `q�zGE����M	�{3��8 m؂��u�5۾�#?R �}�A7-�bz>_���-!��@4��+��N��r�<N� ��zW���P��n�!~0\�q�gϑ[#a��h��h�����P��L�4az�S�7	>
V&�(�f�$��f�ۮ�����f��{SC�7D�8��cx�����֖�&9�s��������2}�V!����t$��G�'�ʐ`e��.�/L3�gz�'.���t�m�WMϣ��R'T��-���	vbLN^Nw`�5R��	"�G}9��aZZ���&{�Cy�÷�#�D��'�A=�G�&���\�(���'a:N<|�%^��pxej�����j�6l��q����_��^�IYC)W���j:��6!��:��`�b;��:�y/$��_J}�E��G� �+R��?0L�ڢFM(����x�f�vuYݰ�>q2WD����c$�Q�����U�d�&���1�5�_c������&����9�5ޛڻ��(F(BM�"��W˒>�/ܲx�=>"�g`�(�J��`{B���y�3��Ja��g�i�i��cQH3jh�Q�990:�O����%�6X���Bf�Tze�*��$M�{�޶I:���S9�=qg$[���ނ�;�F{�������4���E�0�d����a:zl�H`�F�#8�:��0�9�1ltO� }�\]�X�1��S߁�O�xpiovdR>L����sw�e�j?P�m���a����:�͙��������R�����Z�H�s�Z��u.��ku�Z��vp����h-��Bw.������ٚLC�Qd�� b�Q��i�e	VK4I�8�*�C#�J�QK����
O�b4\�I�B���i��b���B�s�x��3N-�b5K%F:�PD��<���-��e�%����D�Ov�����]�}
rU���#n�o�h�ؼU�R�tt�"�:=�Y��Z,R�n�z�th��������_F�@�,�<�,r����`ƈv��v`M��&r�5o���>��`��f�_10H�����5��ڕOW �%����g�A�as���1o�D:F��uf9'�+f�B,�k�8:�1�pv��]���v:1^.��I��x�����H�P>�/��A[�UW�[�[���j)�\7S1�֤�T��mP��}v�V?�ل�*����D�ң��&>�����J�]�;9Or�/�ٓګ*�^��	1�s�t�gx��#&P��@�p$tEѼ�I��Y����d�[P�'Oz�B�0R����H
�x�k+��ԙ�f��qP�Ɍ�~	P	X�v���@���Nbߓ8��JH�_�;��w�ș�����gm�x��]�U�5��2~�tQ�R����É�t������CV�"��8�q��5��|�Ze-Q��	Z�0��@��s��H�"����ڊ5�V����,ɻ-n�):PB�[�����%���kG��{U��T����Qθ���D6�g#�8��z��)��S ~�29��a��Y$���蕨˸a5 ��d�u�;L�:�D���8`.�W�]˪]���8S���Y�϶n4%k���M�w�#cC�����]m������[�L����9P���־��v���_5�Չ�N���dK��QW���C�~���Q���Ae91q[(��9���J3z2.�����.6�k��}�r+#0�1?�`�G�u�Q��a���x9��� �Ew�;n��1xf�o>����ld���ȭJK�[�ۡ�b*�Gh�?��m��?�C A�܅:#) ����Ｅ��r"\#�ђs��3h����:��*�nJ�U}�#�]�6b��ͷ�	����^� ���7&�Hn�\�1A��i�T������͝�0����U��A|ě���L��q_3Hl��]u��"O
��:f���E�g�Q�3�/;�mD>�v�o誈�9p�� ���l���K�y�HD�;���*܄z�ݶ��[�de�d8��bݱ�¨k����֒l��3����vN����a������/U�\ ������]�w2fq�*22WX�(�lz�;�zC��4������I*�J��Z��;�S�ѩ����f>�	qP~Tj\y��a���.�Z
�Eg��&;����;&xΔ,2��l�չ�˅��O��y��o��jX��<����]�4V��i����	���>�sr�?�7�8P�\j����� In
	}�wd��q���L�*�#;����?%���,wG�����M�뿤�1c�������f�N;���I�&�0�,*R�?O-@��~��r����Jb,m��&�V�9O5翟a�; _�ڠ��%)�J�*����[�*7�ي�cӽ��Pg��2G�;b�2�5^h��BI"���f�e#�]�_߳�N�J�z$ʀ�İ�<�j��2�6�Th�i;��
lf{'
(���Cq�W��\���Zڗ��&<h����.Y=�-���\��4۠kZ���?�� �a��`�; cX��cÖ&�s�&?R�,AB��mUP�ʓ���Q~����ܩ4^yL�6�?g������n��=���7�~�G�X1f본S��q�TJ��������[��n��A�k��ׁ猭�I/�+�ݘ�m�?Yɳq�N���fwعs�h�g2�3>�"���;蜅���k��P��T��L�Y�m+��k�1<UE^�#ωF6���0���Q�"����4�V�F��0J4���-I��]�)�Co���j:�����D���xr�k<fV��!I�w�!�;�������.�W���.Å,Zש�k��=��x[��sz#�9�������hw����-��3�G���_�����/J�)q�;�E8��+ɩ��n�}V��p�
��8O�t�B�_=����k0��q�nTߜݒq��`=�z�P��+x�iV��Λbt:`�����@���o'����D��e,ЄT�'��κ�~��g�f`�S*X�w�ossA�:��
�й�4��?b�{T�X�Q�-;�i��p���"��U8]�H'$�-��V�\1�x�N�Xhd!���n�(ՋF��~�j;Yv*���oq%���oA>)���g�&9"�����PC��Rp���C����n�q[��RǞjM����b\��lE���d�\�6�頓����6"��k���S��E*�!�O��|9(b�� ��	�D���vwTH]y�YT~�8�j���͌7���V~j[�a�6ʻ͎��L޼8,�y�8!9g����C�­[д�����̑"���@̠A�D���|��-��I�M3��L/f�I����͵�u��
�T�Q{��O���'�	�E�5�z�qA�\��a`p�&�-r5dv��\6H`��B��)�.>�-+["�4i_6}�A^��L5�~�7lð��p��`������w~u��^�����T����h���"�}�`�E�7�Y��*�����(@�U!X8��E�6�r�sX��aTzBHA��_&,��^ɓtP�>�?�V�[��y;��M9�Q�Z���h1��D�[��$o/+4�F����u9��<E��MO+C���