XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����~ǜ��%	oJ ��0��*�e�5ٷr��XO��"�M��8O��G�,�����(�����{..���Y9�z��mng�Z<��q�������;���ޭ2,<���)�q~$)�\�q\�^R�O6q&�w��(q}�:�~l��o��{�I�����ܞ0��h�U��ƌ��������g �c��vC�__��r\i�u�./j�@J�����)Ryx8��q͛Ӫ)/��mMu�r����i���.������y�MȉA�(p��8π-���Z�Ɗ� �ݶ���,��j0���J� ��(������ �q7RD8�k�@��C��m~�4�)X7����3B�6���u�f�v���4�l���PNc�T:!��b�z�Y�\}�8�c�E{�r�������K���U<8��0D�M%C�ճcH"$Q���Xu�m$� ��L�z����fz�/I�	ȁA\�F,���u��Ԣ���Ҷؙ��BV�D=2O��iE�Ѡ�]5+���W�Z?���;+��ǚ�ev� �oqx9T�����N��(���T���9��d�Hӓʗ�~_
�Fo�wiUTX�4�s>m�ǯ�k�7eV�� ٶ	ma�L/x"Kq��=��U]ڇaw@O����
ms!�he����~O��6i����k ������R�~EN[��q�y��DC&��C��ϫ}5�v.��G�+�|�.Q"2�M#'�O��r�I��}�10�g�C��*��(��-�p�v�XlxVHYEB    5866    1100����5S^6^��H�=�Gy��~�R�oQ�|ܟK9�(��]��#�6�r����s< ������jÕ��7�F�Gs���X�n�"$�����U�*�fj߆���ۅ��}z�||�_B����������=}�3��$Kr��T��8�L�y����Z�[�Z~+�v�8��&/v4S�7˄�x�u��q8Aۣjz���118�R��"SNK?_�����^�E֝�
����.Nz1�Tq�3�\ǅ����I�_�n`2��r�F7��,5,�����6$�UÎǰ�Et��=?��]̊�VeM�P��W����@hN	';YZ�D��'c��Q����r�3Џ�C9�믐4D��T�f����ɴ�lI��XX>�2� ��$6R�>�_]�VP�Ll��TM��`�3S��>~K��PqiU�0�!��<U�s%��X1X��~1�Ϩ/R��0&���9;%�C�!�'���h�x�mB=� A77�Ȳ��7��Ҿ��L�B*��_��5�tj;bW(�����'*R���7�G���~�s�X#��L��J�Kf/LW�uY:�Kf�x��Ls��(t���D�ˁŢn�f<h� ��^����h$�Q��5-�� (������͒�k���X^ԭiķ	���JW��w�t&�P�;�m������C�A�����MEz�W���j����N��BA|�r�Z�>�H3gB8uzrU�u��C��D�c�hX�F��������-�a�z�G�,�
b�>�Hl���&��Aac6wf��S�{���/� �֍�bf�T視P/4y6�'��H,!��x�ӃhiΜ��� 
�-���R<=�䫙2�s)>=��%�v�kCq�h{ȲJ�v�j롧`ė��98�^"���$��(;��܉x���kY�&E���)ՠ��CdN�rj>僎�� ���=��٧S#=˳-l�$j��kP5�?�խ�N�z�X^��4=�y{�D��y�*���-Qh!��Pdf�i�/X�o����k��<XcD�]��P�vg��UJ��
���Tࡵ)YS��b�x��@aS>��9[��@t�K�>�;����Ǌ�6gُN�XĦ����%{K��`��@tؕT$�'�2��R/�q��\�	v�#�x3���:?�YA��+�u����w�ڮZ��L:s(�J@X\c$��s�l��b��(�-u��,��t<S����O+d}!|�j�v����snx�/
�/�T��vòRG;�e ��p�M�s�Ͳ^34{�8�I�D5t��9��la,w�=2�j�,�e��x2�b���n4�`��|�#2�Fk��򶣨+dl<S�Q=�ۭ%�����$���H�h�}���ѷ��D\२R�C�0���1�Vd�p�;�Ze�Q����D�i#!�-�	��dU��Ͳ�N1����C `�*[��\�7��ySR#ZG��/�U?�@�SraqT����C�F���IA���)�P(�Δ���8~��x�ƹ%�5i<�Td߆g��op�q���8r�k�΋y�>o�����J[��bWQ���i�����#J��A&M�:�W�7.�y���G��y��}G�����BD�u@���N���`�8�Y���w�����7�|�kʴV%ֲ���"����P� Z1����2���j�m2�\���k�vxt�ȁ<s�*(�1��.,,�����E����a=b���osR�M�5�L࿠�I�;W<���?sϡ��j�Q��\p9���c2�uo$o�-z��T�	��-��߇��dб]eK,X�����h�%�~`��XA�-��Bu�1$�Wߎ�B7��-S��g��Y���J`��(��J`�.N;�d7���9 0��N��:���ˮ�"3X�s{���O>ÚVN�V`�i���>��n|�#��o�
sL"�w��Z~��A�~Rb�N���[�%e�2KΕ�u<[�H��вvU���_�ǆ��Y��V�'
�*��~}�Z�4p�@E�BS�u�L��z��Hڠ�0ݶ��(��d"Q��ᕁ^���2���aqX#���l栜}�;Ǝ)&�u����������IK�%7�)���5`����eL�$#��|Ϸ^A���/;�HIVC4��|�r��ȭ䦮�
?�x��+��%�"x� -�R+���:5i%�k�q-��2	e^pWp߳� ��#��E���p����d�i(�����"�&����Ŷ�Ӫ���jd1hf%0�4�!eW4�ʘ�)d�v4�;[�Qí���3Vϼ�R���þ��n{��d-���,��MNP��|9�m�[�q��K�g��j�)Q�(~n��u�Z"	�->wi�ԑ�P�R�\\BBnBb�-T����V���l�z���(� �t3�D�O�5�}�Β��@G\���`��0J�A�ϵ|.�l����X�uB�i���`��.�	����N������̅m���0\VR�o ��!0Ff���Sq�������йvKR�{�����c|%�1��.���"f"�,�TАY�y��*�bQ(]?����0��ވ%2���-o�f����(��4թM=�{�N��3��`�Q�Fq�|��^��=�@݅��:�c�1��1z������*�'��y�^H*�E�W�ل��$J��#2���h����AD����x�)�SLx�_�XS��F�:,ylM�X/�uL�e��<��1�k��i�8����S���\�#^���ԓO�I�[�J��W�rD����T
�����
0�]���8ShE�%%C�F0zF� =�����e�BvڭJ�=����y�POdpm3����2|"Q��rԹ&����S2|��!��������l����b
��/�<X}\9$}}��~�c>�%���	\���L�Y��O�g(wtS>�Xź�[hs��:|�U���%�CW��5�| e��nF���E��a����JIu�]fWВ�1���3c�.H���T��U�%H��5R��/�O<:�Aw@sOO���6���]�욬��Biԥ�9�X��Mn����唪3�"s�sy�-ҩ&����s4%���� æU>���#�Jv-K�y��by�,�(��j��"ҷ��y�\n�:L~�xa�1����"ّ��}d��x�:��y�q��7������Z�L�g�Ӑ���!Ӷ�+�hJzj���'�l�IQ��2�oC�������Q�ێ1B&O���sԝ
�[�p~\�ʎ�w]$�yqjt9��P��ܰ$��c�-$�E�X_�`u�d�4t{�j+M8�'n�r������� CJ?�z�6�j+��fJ��������T$l�$��M�3_
7K��?�h��H�ىt��2!D���A���v��k�i�g�I⇮H�LHh>\��ʹ��5�wzW)�U�9�.��G�V"D���el;̣�C(���<)u�Vm7���*г23�T�a�]�! FQ8��.��
 6����_�߹�������0a�̯��~�����il���
#�ZD"�����n���DAe�QN�Ҭ�;Z�Μm���AȎ��
�T����FwT^��K�(�Z)l�^�f�~kX���k�"f�W����ET��J"{�y#���?����e�[g��{��SsE��$
����̤���9�vӤTsX|�k�v_@ ��$�|O��4g�mT�lSѫ�fNz/"�h�ܑCc3c�]L1�@�<T���&�� "�<���k�02Ǳ�X�AI}�8m�˝
�(�	p��ں${�w�0w��mIF�Otw���t�h
'�8�s�+(D4X@����^�{�yy��U� ��p��UV�+��8�+����Pt����SZ\g�'��8۟�s�]���Q#5BB���7>%[��(/���#��N	�%�B��d�A)r���sf��}>��u���0s� �%g�4m��)�����ޏLQ$������v�Ej{��8
�m���#�Ey"ْ��x��Q[��r������o�!��+��q�|�O0E��}�Ԇ{��^yݦq��@���R���I4R^���Ќdx��%݌7P�Z���13�q���*~K�b�t�{f�۞�E8���%�R��Yo�%��w�DLx�|D�g����w����(��	|���C=��|`�O�������p0�@s�"y����oMgu�gY��\�V�\���Ab�^sr�Z�uOp�e4Cgv�����k�r�w�,��|m�s�S^���mЊH0�'��[���">A.A�1�D8��L������