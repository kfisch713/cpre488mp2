XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}��[�/��&W)��ĳ��RB�v+�|�����j�-gzk� X'��N�^s����ϧ�pN�V_
�FMh�A����7���*b�H6���wOO���5ߪlŷ�չ!V���` *v�b{>8�t�c�XrVd�Wp�e�5P��!jbG�-å�lY]��%B���;ËC32/L��"
��C�r¯O��f��mRr�N������4��b�f����KhNIbX+_��7�\�I���h�s���G��%XYŁ� ���(��H�	�,/j4it�"��,_u��N� �x�<s�At�����.7e����j���
A��=tC�o����Y5R�m��!ʤmHIM[��&S
'`�|�i7�i�*b2xcQ}Ŷ�����"��j�<2N�A���1�ϥ�7ys��f����ݥ�7��!m�xՇ����zr��d<��(�&����3	�/
��~����u��5�l'�����;�� J:�9�4��vt���.߄)�9XFx|���YD�v+��h�����W4SXhA�_<�Q	3>I�m=�v�!ª��!�7�k�M�?
�S����h��3[uz�7{���}�>\8�0����^��B6ʐ��|�������DD����Bk���Gp(IJ�b�^I�4�ꡱ˥ۃ�#����2���=�`�cANy^�[��:x������&�J�u9�����m��d9���-�a8+�4ѝ��X�%B���#����:�:לD�y�$����XlxVHYEB    15bf     890��+�o�� nGE��0qI P
A��|T����zG��O�wW�U�����k���Sq)� I�S��OP3��d�X�L`Q��~d%�q��:-�G����{�8�9=`ɛ�� ��;�
�v�d��Ľ˻�v�� ��T��}dE����D ^���S����NҤJ��V{$hu-���}�?;B(ܿ��Z�!�z��,�\�g�a<�O�8*���;��Y�[�q��8��3Ɖ�U�&�����B�`���Fx�˓t�V�h�r�̰!����\�l�,&�?/�t���7�ϱ�m�%�����k���9W�UL|����i}��
9	����z�~*���7Qb魦��Q8�Fi3"!�c,��d�`��J2^���?#H����Ϳ(��j�:s.�zϚ����҄,g��/�e����i�6��"������6��t��o~�d~�h�^�I�5}{ �a�mݝ{��P��fDi@3��zq(�3����g���mpnXtP����E.����i඲��vs�?�����ܕ��%ަ������8Ͱ�V�vw�؛�Ѕ���W*�u �y�Q� |A.��2-�[y�~b�[C?_��ͯ��"�vv��U&�TDk�Y�o�p��~���̈�;94�J��-����J���n����ذ�;.��	4�j���L6ݍC���LSB��d~R����1 �A�X	s
�:�S�� ��5f;��j�Bo����b�G�p4�F�B-�!�-Ns�/aR";Ѕ&��C��� ���^��,^��gD6x��J9,�X�-��a������btb-��w@������_�ۨr�����[��Uz�����nh�)�C+�{����U�L�I�G�X����^��f��U�R^���X���6��q��ŷ�Jx��!l�����X�$v#�QhW�~ä�����x6U��Y�X<�G�w"����c�:�k%�̴60������8/Y�U"�N$��N��6���j��^�$�?C���b�g���曗Hq�&ލ0V��q�p��O�
�(E!y� GL!f��W��/7Á�ь�@;\�����4Z�/XΈ�5��/���kZ;	�� 2q��UU��*1���i��� �(�ǫԠq��a��C�[��gDҨ:����7ε��b�N+� ��ax`z#�:ɸ���TF���C=U��9��5%ΝV�P&�J��b�����،H�j��V@��-�1s�RIeg�=\���<��OS�-	Q��
>D3� E�P|��j���lͅ���� ��T\�����iVgs�M㞐N��o'z�d�
���݉ �jP��[N�Y3ÕjZ�<]۱�]0�1�9����˽�P�7x+-o\���L5����%!��/�K���D���<{�^F��G�8k��:{�_�r�����Q�΢P3
�ol�c�0�� ����@���.Oz�Av�s��>ce�9�w{1o������"�顫f=)��� �6TY��J��b��FA�6��v������P�O��N6����z��yM��3%Q3��a��(5.������s6�v��e
�>��W��*�We��-���inh��/�ByV�;�y3��~\}6}{�5r�W!��b%jd�+��Nߘ�e�kq@�Q�J����"�ܤV���-U�u ��r�y_f����rzH����3\7�Sp�$�4��MfD`���Q����d�?��%r�^��?"���朌x�#�1$�� ���l��WK{������H�ǖ�2kl�kj~I	��,a�@��A�#�bR?[y�2���݉w]�+PS�9]�2e��>A$�U�(�gt2C-
jp��u�,a��&�Y�u3d=�� *�>�-�e���f����OSjq,����A�������'�nw�΁ؽ�gk����$q&��s�(n�W׸4l]���J�J������\���&�U+ms�dX�pB�P<Hʛ�z�9�B���a.nB$�@���OFx�o �<uXW���n#!�
 q��&b��;kx�����T�O&�Ӳ��E�����
������8�7��h��ڔH�`T��3=yK#��H4�T�hg!NK�]�$��~@�G�����#Ļr-����P��.�F��r�'��s�raU`