XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0�N��y�`������#{ސ��k�ޝULKG�6����Q�9έ�mkFc<#`��|���yP%���a��u��C�Ω����#v��18�Ao^yV�)�e�����\8�<�@XV(8_ds���Wi����KC����x�g �u��y2�Ec��c��a��a���a�'ϡ��$�M����s����6	�l�Y�G"&%S�{���ql��������1�~ )rVa8��%_�Ŗ��3�ДH���X��O;�N���We���U��bş����������ܶ&;�ϧ�H�4�z<���u$F6����u66ω�G� �^A�@#N���CaIf��OBy�Cy�����F\]s�WTf������V�O^����,ۡpy��XR��^�2m�55¬kc<[ @�uD1�	鮪��$�����U}A&D^�c:�-�t7��:��˶k��6����&��\��D[�̄֨jQ�FpX�5����Z'\�y]B#�4`���Wf�x���6��0��H��&����B0��ahe�u
R|�%�ey�Ж��m~^�e�G(�X����5=�[t�)\L��)���K���#�_գ��څ?���C��9�l����1?Um�(b��pK>
��u:�<�NT9�'d\�R���wق��͞��5���mNe�H0Z��P���*l�	�W� G�%X���y���f�.�n�!Ï���I��o���fF�Q�B���;��WE���!���4Bٛ�
k� �H�����k�U2�XlxVHYEB    da59    2e30	<xv��� �b9�23雵��m���HuA��@ 9�^/�����f^Jŏb��Ԍ�47}3�RgF�����t�5&��eh� ��r*�N8>q�+7)�BQ�4�Z>_�}lz���e}���5���s��Ƕ�eN5.U�������O�:��Mn�(.c��x���wr�OML�R�a��߀�0=:�+~��f�4�A��I,���Z;"�bu+�M_��z|0$�x��'Lo�B��B�/)X��b3�g�l�>Y!��Զ�9ʃz�����B����Ls��'���h��8kYDp�ub͕��ܓ��}��!�P�Yg�C�4''*O5e�yiRs����hcO�?��NI�^X��
�����/V��p/��>��>��Xѐ64���-�xMHY��|2�"�����d��|DN�Ip/4�1��L�/�wRWǡ��Q��OF)d�E֥�U,&�E�C��$�Zm�����l栓�*ޫƺ��aJʓf�Z7��C�R,�[H��F�+���_��g���]}_�$�I�dd���`�y��,�ŮA��))Ʀ*�n�����S���?��jĮX7k�c��o�1K|ܗ+�T�*c>)���>\��(�~��zw��v��'�z��z����o���JI!Y̘.�7Z�������>�5���EM(�u�ֺ�����ܞPp����l����5�Fg��0,".��6�ߥ��i���bh�2�4��_�Y0�/�F���1�6�W���~G�̪wV�M� Z�!(�Q�>����B�Ҹs�v��kc��[��i��o�`qP�;�D "��D�5X���^���vP��n���w�ˇ��x��neH3���T8+ܪ�F����z�˙
�Ya���BH_m��T�xA������<4�� �����#���>]��	%����]{��s1���K.ۊ�ա3ZI4���=�������+���P�1[�H�g5`�dv��D��w��'{�$��6++�c�k)^�A�4?A'�
8s<�xG�s2�?�v�	��9DI�L�w#��4�l���
�N�Y�ٿ%_�Aɲ6�?0�1'�.>0U���78P&!��?�c��#�C����HXX|��&I��ެ˼y����v�Bi�](7R�@��a��T��w?��pm��D�:,��S�
�'�o��oz�E���Y-�"��;��V�u0$! �8a�pp���|3vσ����yPr�/�*�zn󛮒��A�f�,��8V�p��t��:�uQ���C��۵8���&~+\�J��F_�υ���P�>p���4Tջ�7�j��)���2W��*����8I����vB�7	�C�T!����7c�h��䆃~&�9Ab	��>x�B���>�X�RjJ�������,dw��Qt�(�,?�r�n��}ؙ��jbJ��R�����-�A'�#o�A����^~���Ld�s&r�������VE����g��.Z�\ٯ�Db�4Cq��fr�b|gy�3\݅���F-�(@y\�d����H�����pm��}��h�<4p-g^[���,��EKH��0�e�H!^dѷ���Rw�~
Voh"��K������;�ť����s'e�Ϙ�"��3C��������cs�S�I �:U�/uDN5��4�t3�w�@�� O.��,��pd��&�o鐦���>J�Q�m��2��&�B���*1�H5Rk~5�U��d��|���-qaQ�Ƭ��+����<'I�U���ͭ�
�*�%K�y�tVV#Fq�U]��2�Q�Y�uQ�����1���7?YMI�V�
�b����M �uz8�b�E �j&s��7�N*~�,�y,A7J�Lu�xO����.�Ŕٓ�Qm�D�y ��oU���H���~�µ�S�FŔ��N�d�W�LH2��k:b�iҎ��<G�I⿽�<$;$d� @� n��oI���|6�F�;a(��?����"��Xa�3'V���dGW��ݳ�,2a̔:��V,�ԃ��5���N@��1Ъ����*<�8!��a�a��~˳��@r����V2���*(c���X_����u�Y�F��q����b�5�3J�'��(3��oL(l�%+Y��<��(������.��(Tr0d�V�D)*�>�8�����<�#��!�����=����~�t�R���	�غF-d�r��1ԝ��U����KC��Y��R��s�{���P�B�$N�sQf�IAg�sQ���h��TA�������G��\pB�}2�3���e�</3V�
��w���A0`�(�<.�;�ߐ?-�zT��MY7��0��^Q��)���yY�@$����[�rdeҰ����d��:ɉ6���:�ֹz��ۈB0Y'c7�8��J�kcj�N��S���������X�ZD�9��N�D@�ܭ�L��̅��
�f�HP~�ez�;�:��.��Z�Lu�����&�L3��J���uGԋ2�[��G�U�M�t.��=���=>9���&Y��h���>]�ؑk�-���Y���׭e/�7�C!-��r�0'Z8).��&�|}=��DG]��jq�k���Iԑ_D��Wڡ{���%�v��	������Y4�`3x����zVh��iG�	t4&�n��@���?��`%�P��~��i2/�A_��+�lP6dh�4�V�H�y�.�вT�/��p�!���`R
�jFPKf���pQ�T�������L��7(%n���J$z(�{�����d�&L靕,���^�e>JbS4Qa״���\?���=qJƟ�ތ�MIc8�G��)1CC�s	Lo��!�0�D�q�=������~��"s���s�Bu�[QF���<��t��������A�J/�'-H�lh�#�Y/��?�O
^mI���=)�&���Lz���?��� ܥ���V������W�Fɶ(O���Pp���(�T>��!�8(ɳ-T>EP��[;��T$��oxNެ`�[+p������Vz���s9�EXEH;�?S��h>`��,4[�*�W�K�7��͒�ü��(j��h��4��>��ti]���Df3S�0_���W4��9aK�1��A�3�K�ǲ¿�#O���J�h��kF�`2�_ug �YS6G�w`B��.�����~��>���i���^N��Z��"^����z�g)JkD�p�����v�е̵NM�M/y"֎�2¶@kT��r�{�!�3<������/rO�%�}�\qAJ�~�+��2Y*�H�Px8�D�e���o=��lq��Fۦ1Je��|�Zpt�����G=��g�h��az���C�S��*�V2�;�⻘h�0��dX��lD�<j��B�Br�Bf-1���!�</����%
����Q&S�E��1'μMk@��#��:ޣ�������I��e�ns��T2�2w�j��+����j|�̃�\�c!@�mVvG-k0�#��C��~��<V`-���"���!Č'5.J��W�\
����h�J1�#3]?�E���5z-�Ԛ�d��cO��S��fY��DN>t��7�7�z��I+FMh�mqg�Tz�vDa�B�~�	\rrE�e��,E��~�;\&��eW�O�V̅!��ӗ��.�SI`o�r����l.t)�=jDAb�'����	�ʩg�}v�]�3�9F��㶛�.hΧ��Z�,��~�ц�0(�������r����y����T�nOfw�qU�~���݇��#�D����iDX3�F�8L������;�̍�(�y���,��/81йoo���T[�p3R�j/PIT�cRë��R���j2{_��]Ȋ�о�Wm:��O��M�%MsX�Pp�/z��{��QY#}�P-W���ڲ�88����"��OM��m�����v�J�d����=|q�Q��pf)�҄���&'1�rO2�]�^�BR���G�����->e��1��o��p<SA7��͞�QV�(�F�f�fFb�݊o� N,�e �v�ϻZ��vq��`FjD�xu��.n����2 wjS7�b��O0��
c����º}n����-����;��ֱ��7/� }�]��Н�<`5�T5�`o6(��Xz�#��!���9��r��վ|����od�!:�#��j�)���elKY�%?��"4�M�����b��q�`����bV���cF-V���� �S��	V=�F��g�v�i(�B~��Ъ|:�@��@q[��vF�W�I��	=>�gF=�#�
��Y=�P��P�K��f�H
��8��k��������.Ct�"5�e�G�I4��>���c�0�{S��]��0x�,�0��&I��3�UF"q����Wq�-�S�Č��Is�����9��8����Y:��g��=���HU�H:�s��]X�������}��C�~�r��69��گm�z�*L���ۈ/'-� �R�!����;V6My�6tz�w_��o��;׌��I{Ȑ�Ŏcr����ɡ��C�9�8|絠�����J.7�q����k,T�/�}�)��=����Ȉ�3Y*��,4��h��9��ga�ɘ���)�">j=JAg#��A&9�;=��`�wo+�?�99S�%Dnވg�CI���X��\2Ym��$��:�`��1�� ��d��7���#�+$K��2-L��C!�zPj^B��< (�ehZmk�(�Vn��&�h��5�)��HYgc�W����יA�2[���i�"����л���%�� ��K���A�C�HN���M���\�v0�
�fY���$��v��!��\�	^H][�ɌL��������'Vj�2QSm�r���C瓽+�HuNJ��������[�W�%eË���æ��,�e��7.@7A��2?Mb�G!�<�sq�k"�tf ���ϸ@�~B�ʰ�cC���t��/�4,	�]`e,��Z+�zY�Z��z�MU�	3����P�5��x�T&��7Նz��Ua��~���:L9L�eRDQjE��Te�����GC�gV8��[Mޯ�au��"<�Ė'j�S���?mMф9)8ԉ<�^���d��X�靭�&y��p��}tN����
.�E?�U�ߤ~�<�ՔP/M�eQ�Q�"��ί�؜�5-�Q���Ū��h��O�����O���B�bw�ݴ��� ����Fj�m5l���Z�#qle%��`�>����6��Ae���fڹ�"SP�T/��QF�g�!P�q�t��4�(��D�HI���'�4���0hV$L���6�|t�}n^��eK��7�#y�œ�~���5P���K�6>pg!uca���:����p8-�[4��6�O7U�?�ddK��1���9��a*��*2_��������W���Ǘz����OG9����f^���P�
�A�@�oS��s9x�e3���u#��$� ��TS���Ц��{�8�f����Џ�2X	�bl�k��!�|v(�v�?���>��\���abER� � f�M�?˸���@&!��-*���>A|h�~^���â���?��RMA��$|:����;�f�Z�z}v�	�#�,���YL6�-�F�s'M@�Py�X�)Sp�����3 0x`���&oA'��a��~K�~P����$0�p>
W.�R��W���Zhr���].�ۙ����OL��m��4��D`���@�:�1�WbΦ�u�o��\Yơ���hk58�
7��[�- �{5T�f�9ݣD4ꮟ =ލ�P�t8�Cu�ʌ�D��ӿm����7].������t3�Ӕ	���M{ځ<�?�3���b�m�}��%�� G�p-� `ETOb��;2`��46��[@l�Q�G?�)}������[�P"Pl���[�^|��L��@��/={є�Z�0��3���vԠ,=sމ2�������T��r?��&���C0�CR8l&2�d���9�!k�Gd%]C�C��wX3�8��U�.$���"lQJ�ֻ�=~uiA��b�oA�|0���uW=��ab��	W߭�Mi�:X�ϒ���Q�t��r����H�1���]b=���j��-�C�b >@���0��ʆ��Ġ���X�VK�m�'R,�Ű��wS Y����x���A�np1Rx��g-4�����r,x�-�G<���ȰŻ�{��z��*��^�ּ���9nVm�m������w�]�8&�ֲI����lv�kh����ǟ����T̠�N`���ڊ��|k��J��K�i��ܴO�Ɓ��֛���3��@��~��).��F�#��q��K)����ҢB�_d�X�#� ((��\w��tQ]�9o�X�釾0�@T<kb��z�U�B.E�Hȗ����c5d��5��含������?X����|vE���k�fq��U��F)�T�k�;\�����p'@�z��t�Jұ]Ƙ��Z^�s	I8��hA#��kүrnK�y1�8y�vJ28�G�d��%`n�8P�R��F��db;�̵���AL`�w/�2GA�3�#�c�v:���P���a�^�>K�l�)1���8.X��f5\��ˋ�k枦���zdD�$��[�4p;�c�s׹T����.�;��E9p���"��T9@��U�G�w�-�c�Y=g�3��kGM�$��4�����s�kJ,	|��V"1��q�t3�m�[i�������.���̼����A_[~#��zO�m�s�%}9��zv�vT��@H���rkR�;�u�c|�&��1�j���W������F�[�X������o#g���������-�*1e�ڮ��*�qCW��X��>�?�u_#�R ?{)pmmy\z8�ɵ+%�Ǘ�C(��C�����+U��[M�+`�su#`3Pj��y;��Q��Y}����?h\W��jH���~>�i�
�Zy}����C���B�)��qw�m+�ֲ��v�����u�x�m}���BƞK�	WzS�Z-���%���5�0�>GԵ.��}SP7�>���gtz�b"��}|Fn��e�IV;:j�߷隿�Vfm�l���u��7��rC�@v�b��������}|��%�Z��	 >'�E晇�.�&�.��4�Z�2;�$q�+��U����*�:�g$S��T�nB{�hrft)C���a��l����!�aZ3,Y9#��&$��5��(2X���p{Q���|}�2��ZK���'���h"h��E�AExG#n��O�f�����z��$�x�p5���<���Hmzug�P�����Hk�5��[}��c�ʁ�(�k��V�z4	e�'Z)�UQUt.�o%j�n�?&O��0���c�H�wD;N��B���k�Q16��&��#0��$���0�8.+)�Ua��Z��ߐ�6m(q��~��W�8�%d��#�,�ș�r�/��M�߸���!��]� [RY!>�Ɣ�����%�
jv�Pe*<�D�l�:v��e�O0B�v�^��F[����2��OO�����%k��g����8=������&@�DMX�o�ntD3������N��C�a�4G��8���ё���Y����$��Qn��������'���l[��[o̎��L��R��߹!�N��:�7���*a�z���N^y�s����>���oY��qSc��3w�E�V���B�a[�K�z5T�q�6���y�����[X�Ec����-�k�PZ���(�3�O7g���}EW�����
c�����i��aY.�ܪxĤ��P�G��ՍieNd��t0h�C��D��i����j�_W��h�2~/�M��/�i`eYr��h)5D������ؓ#�,,MC��]�a��;�N�_o��>c6���|_��ET�vgL��,�5��e��sǍ#���� }x��۠Lm~ˍ�x�'���G)�N��F�8���5T�a��fe�&b_����n3�]AN�6���:���WzH�ܠ��\�SfP��Dpl؛� �$�%J�;��=����� An�L��?�5�M��n�/��w�+�����~Wb�@�(WZpF�����cg�7���BA��m�&��X]IS!�U�k�?�%��� 0h�O0�7�sG)_,���JYs;���X�	���Qr�����y�X=���Q�x����N4�[�S�d��HQR��_e�N�LZ�ѦC�o��/��H:F�[ߥ���m���zI�N�� ��Mq�����h�#�V�'�8ktk�-����kK1$־:��+��ȱ`mY���pzmc �o^3v��	r-M��.��ov0��-k� �6D%���Ϻ2M)9�>�e��eK��!��-
�s�u���X�Ǩ:>��k��#�) D/l�7�Sw�___�35�bhX-�܃U�Ï�aW�T������4Ym�-T:އT������xT~��-��Ƒ5<�p�J1"��D~��J+V:�e��~P�f��VP0�ᾛ��TEn;����ʭ)�����ﹽB�p�HTx'���!y�nĹ @DLp�s?Y�-=����r���g@w��R|	3)�Ug��!
J�#��J�lvVaK�-IZ�쐰�	��F$H�<?*g�20����c�������EŠ��74U�9�6�6�/����1Dr_3!lh����tX�B��'�������v�� ��Q�����;�u�u%]���y��y
��}P%�V)��q_� ��^���CtP����7��{����wYjg�:��%������ׯ��D/}�r�x�s��� 6s6�zwr�=LP��e��t.��Ն��[�[=xZR`�ao�'���|��_��_�uP�+������H��JЦ��>���[)�Q�yn���R�e��]��,-V���rX��T	�3P)\��@4S�u�#�"(S7P�� G����h��g�����#Td����d�~ֿ�����˦��3�	%L�m�s��D�{zp8�^��K��>/���SčR����?;��?wm�Q��؃F��Z��
|Y�5/$WF��.��' �o�&ϻ����-ԍ��D����d���Zʃ�"|]��E�x0�Evz�����h~(�^}��ݝ������<gL*�D�cx�U<�m�a�|��e��DJ�Ğ��u�?	�TbgV��������9k���]9��5�h�L��6�U}@Q��ț=�kP1�+���P}�U�G.���uМ��̺����i>��U2���P]�� ��菶$]�'���m/Y���y	�&^�~�{0��d�w��K�}G�Q ����:�#A����J?S�_���̌�Z=*�c��*I6a�y0iA���Jir�OU�������2D�(Kz�i�l�P!<�ރ�hiU��xpX�)�ڰ�im�W�ϣ.6�h����	���5�3��l�8���O�Ǘ�H����O���?U��~����n�'#�v��A�p��r�������4�kM��Q�|I�B�>�\�C�u�#T�0����b�G'K8�}bqT��$�"w�����=�a�<o�=�P#ϻ`���$��k���?f.Yfu&��-4�7����wa���Dm�.m'�d.�ER��l�%d�A�-X�
]%6�� J(e����8{��'�i�E���}n�+��ko1�.C.}H�×��[Fqkou�R.l
� |�LoN�P�����O��.W3#*E[G֓�̳u$'
������)T�c�y��4<\4�Z�6KU�*sq�`gei�W�
3P����"�)!._P��oK�m8-#����/ěv�����K�u�{'R�v�n����~UCbl�7p��s,� 7�8����6薭%:���,�M��u��Z��N	Tf3:�̓,�\��[48��Ȩ}��t}u1��t��?vY��^�����ԿKN���x���uQ�{}���z.P^&H�L	��yN:3��ZX�KB��i���X�o���罅�����m�*��.6>�	�htN�x:q�V��ξ\��]v�{��1C��}�-a�.2ݵX�S���	��:W�k��<�SϿ�6�O��m�fq��h�7�0C/C3�`{�bV3��U@��&pIhi(��x�T*��D���<�{��_l�'\"v�x��i�ah���K�&�d����0#!@�1�즅���}�J�s�wc��XQ�Y�.(��=-�n�{V�&��2��N�AeP��D���<������S����s�xp����S��_s(�#$HZ���� v�ƾ�M�+3;Zۻ�z"���,�A�����9��5�P�b�2�W���^ĭf�͒`q� �kl��J�+���W�-�X/�'�V�$Eio�z�0r��D�M������;֘��T1�a��$�~'M���B�V*ơ3�vܕl�5u�]��j�]��z5Fn�h�q���i���Q<[��@�X&>�ZX�
uQ>����f��Lz�Sb���b�kd����������Q$+'`��x	���H�oW�\_Fu��J�CoPB��H7*p�D�g쩌+����T�Vװi�����Ť�V�B8�Źpu0�2D��dY��o,8OI$�=��2��E����Qa�c]����ܤSW����F>� >ۜ���0�iJ��z�(���t�Gi� +���֊5��&d�b���b��	6�X�.����'-6�#G��I|8���l��s�����s��Y�n��\��?%����A?��΋�.-�0^!!ظ�B�Ͱ�-�E׾~���@�W�D�H���@���Xıi���kז��FMD����o��EHlf=Ғ�\��_�Xq�0{`��v���6��������u���+��6v숑VA+4��1�}�^<��eh`�r��+{b��"�:C���8��0��@}���{�~d�ΏD�uۚ=2vmG��+P�,�4 ��4��(��H5t�>ڴ���=�N��~�o�����^�h`��=O�X�4˶t����VZf�v��NJ?{�䟇ԍ�p�@�r ��	F8D�����
֛
`��?����$k��銾0��Hۤ�k�{�^U���^��D��STY0�@�X~ת'⛹�y��g:�ć3��'�[L&��s��#1,y��`$2�O�����A����\�*mH%S��iE"�O�k�F�r�����*��|�r��pe.l���+a�p�s��;a��R��(s��J�Ԇ��"��_�ס�iD๩5�=2Y�[׭�\70Q�Sp
�B�-�R���(�`��'wX"��)�w"@�BＣV�m��V��l襭T}�{�,_�)��e��2*L�h��譁>n��&�F�M�� i9���8�:$j��^��E���.=b��A&���0�(��m~��Hг�����9�h^����	T�`mc�T��_� rCP#N�0=A���i̙�@k[p���X7�e�)�2}�[���� ������i��>"x3�����NsǢ�,��x7ܦ[й˄uL�� i"w����޻��C	�>�'[*�H���e�O�Ts��+M��Ka1��f��]�k���R;��˝4�p�=#�o��ȣ��>k�S��$�5