XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����-�Aߦc�}7��癍B����s&v��P�a���e���t��u��IB���y_U�4%��3AW]�X�
�k��-��/��(�1�p�o����G���d�����-�� �}����|3���jd,��P��&^y�de��̧���4&�+���K�C�pB�{߼R��?Q���+ "8�S���Gz6�?��@�����ՠ�t,qA�1�m�@�����&EpAP�}2o�ªyt���u���vC��� �j����{�Sc��C���xʌA��d�UdG�X��:z��}�^'���e/J�!�����U��GrDp:*Kt �P���.6ze�����w��ɣ��O�RI(:=s�St�i��p�%tkR�s���{��7�p���t3�9�^�ҼDs/�����a&R	7B�J�C"�U7^��ȋ<�p����f�u�[!����ׂkN�Rep�=��j>�JT�O�=[��$4�D0��QO���__�6���8� �H���h�h/����%lc`#J�L���f�X'��,������2#�KL��j���{&��ŎU56�i6v���>Hz���DߔqK>+��(�~�c-,N�-�A)1�p}an��{�h�t�եnzu���:��˟c�
�����0�'���.�XZZ%a�g݆��<O"Is2<����c1S�D��NTtLu@�7�B��S�� FI�U��m�(�� /;�K�(n/��X��C��w|	�)���fNv���N4XlxVHYEB    39de    1170����?1�'��u��w�C����f�PI�*����1@����H��bU�h*��&@IU���>웋P�(��0���Ɠ�=��X��w�q�� iy�KP��6�B�7���RT�_o����mI�hv���X>���Z��T���N��Ծ��4K�a�K~���fu��A���[}J�$�����q��3l���-؃MDz_�Q�?
u�r����d"�4=Ty�7��� 9N���to���
�k
�5��ѻ%��c�n���e����o��h�7m����{�ѯ��L�8�� 酏/�qӻB��!�u��W�ȫ����uJ���$����1?�.a�_O�Qv~�b�FÖ�j�6Jg��Đ�+��o��-[2����b>$a��D�
�Ge�7X��8���E��
I'�A�A�+��K���+�F��Ҥ�gg��j���D�44�d��$0�!�1��9Ҽ�k����a�g� �5�v7�T���1Z���p��Z�
�;y������>"�^�/����'�Ex����۔��"Kq�y�P�m�px&
�5%Wʿ_�jW	e��DD%��Ñ���2�L�X���,��S��rKTs��:�a�/��@�aSxA�A�g�,�����\� 7UU� ���W<"M�G����F(:=�f��mKh�������{ >�c������-�-N����g��H���u݋���g�n�1�$�����DL<�H�Ƕ.{E���Y�Do�A�F��9��1��`؀T�ZV4�vs������hM#ž0S�2!�}�X���J�&�?w><��}x��Y���L&g���&�iڠ�Q�u����i���?�d��+�KCJ����+9���@��
r4c�dG�����w�b&"�$�$?�\��|�wU��s�jˋ�LgIG-���W)`��N�B��A�'���U���᭄@s��z,�Y���x��T~���4EGh,���M#>A��4oH5ܵ��^� Y�~p�z���!F��߱9b�����F������NO/���'k���fU8�=�98��]� �"����f֯�R/v���_�g�4��X�9~���.����W�ky�P�k�����d���ӲO�Py�`��l'Qx�>��t��]N�H-,_�Q;�??u���ڣ�
�qfZN����e�*Ɗ���I�s�ݣ�\U�v�pq�����3�@��3�CF�qniڗ&,��v��Qe_���·�t�����J�T�z��+��,�Yͯ�6�&5�L/���tlU77�]�îD� �����(:�(�!Z�~h��mx��QȶC��0�x�)+���EƙސW~�e���Ɠ$�vn�p6EJ�n��A���Hm_Wc�b.Q�A�zdm\�qW�u�����"sjy����@׹����q��,jqebȱ��䋜�/�%����r #���W-}S�H��>|U6�~��(�&�X�
)w�_CM�m��eP!e�!cm�������w	�c���b�ߑ��r��wk�|g;�[R�*���lb̼�e����E�1L�ZeT��^�7fՇ�r�����(��U��G�	M���=��$�t?7����=�ݺf��:�� a��M�s�VK��$�#Ð����0>k#�������\�x�k�t(�l�ۊs��w���P��U��I�v�J��:
v'	�Ͽ!Nٌ�'�3�4?��_Z��Ul#�S�B�tIC��˸����K,{�~?S�)�,���"�����ĎX��AP��q۷�H��4u�5a���i���o#�C<u
\�>6�FP�C,U����ݣ\�<�i/	1�e���P�(�.N/R��7Mk���_�hT3�We�$$��y���@$'�'pȇ|���w��'z<Q���:���^eâ-�p@�K��� L��I��H���t)
G�+���̤ 
����.?b��]C`}���h�E�ё��8��'��N�B�@�����V)kb��8��������z��k�9�1a�L-/[��)��7yu� (�ku���M$7P�'ȋ�,�F�+.�n
����f1����wCZ�ԒS$��ү�PI� ���33QI]d5)O���U�k6�K�B�l��*@b�nZ������zL ��K8�~R 3�X��l�ޛ�'��}��H�E{�� 2�z�D&��@Ő7��$T��a8�T��ͮը<�q��\3���
:-��a��e�u��z|	������������x��l��]O>�����%'PΉ�lNA��k[P����:��x���]o}��s�g��آ��/�����R�C�b�
f�γ���>��*\S�}���Z��4�k��t7Us�Q�g�����]#�?�O��)���R�0�##����ï4	y	a^�	�\�?U.N��zs���&�h���(I�.nͮGB�IJx���VB�g`�C�1ؓ�Հ�˖v6����PhkޑU�xv>BZ*OQ��y�^����ژhǩ�u���5��K�Myy\�a�L�ݵ�RhM9�� �Y���^E�;���4�E�e��1�c�!�%��v̱l7�W�9�}���K��,���iU����+o�ɯc*�lƂY-��r�V���F��	?/�+�f::Gӹj��tƹڼ;��^�S�egXM�Ǣ�ɼ��}����DZ	�c���X���W;/
�����E�	@x�!�{�ϭ���[!3�C�56M�Y�#CD�G
�����*.��r��N	�Ҋ��Y�=�R�	��(��̎���ZF���Sd����|��Je�_\�2��R�2r��KC���#Pz�q�9�̊����N�H�[Z�
[�$U��D����HhW���(��=U��K�$\�h��H�ң��qzE]J�8��� �UZҷ'����(���|@���e���y���e�k�0ͤ���Q
�:����;���Qc(ZE�-pZ
z�p�T!�ԟUv�@ȁ3;/�O��VLL�s&��2�V�X��64zW^��B��U��>����}m����fQI�R��^�9Gzq"/Ja����d�J�������^F)�Y
�ۦ�Q!����'b�A������	�}���U�9�Ki������E��<�c�B)�=Y��E�tߵA>����0���L-�7v7�A�@�`�-�mjך������(�*<�s�k��!����5���:E�
��3�0�յKM~L�M�1�ܲ%��2�w6����E�˽a��v�����
�� [�ZPD����YQ�'���[\�g~M���F�+���P�X 8m��`�z�w7��x��4�V]�*�ˑN�p�Q�}'��Z�hu�&�4�D�m�^áψO߇�-�So�q�!GM��EN6p|c�!A��2�\)|.�ҹ����А�PL2��Ý�ą��MF�U :��A��&��a5�C���i

��M��)�\G];����D�2��Yd��R�8�?���N���J�\;X�/�,��Ϛ���ОX���h�a�����ha�w���o��"�cX78 �5]�
m�����Ux�����i�nX�u�rŌ����i4�)�K./y	���77Kx�m��l���\�CE a��<��wnD�@�r�]��Kq��x��) �;����xz;�t�j��EI���Nu��tL�! �-W��n�G�6||�k�I�
�ϳ�ہ�'Rf��(����v�G�>^39'�#�g�SS�����A^���P`������T�4Y��O�?j�ko�_ƶ�{�	�NX��]�}�s�PLޏ��s�b(L�]�G ��aZ�WS]�H|#�y�	�������'��3�U���꾋���(��QȖ?QG���բ���'G�
oT��+)\B����u=���dAƄ�� �����j����קVCd3�E����p�_!E8>*0�=�#4i@s�v���7�y����e��֦)M���ԯl��t^&�U@�~�G4%	���J�#U�/�^��_Mԧ%���Ӟ���zx`�^GE��Kޭ�F�KL&����e��ટ�i���q� k M�N0��\�I���2�S���##�N�'�׼I\(Q;�/ei��^����m��x(iNݶ��d掊�:�����������誨�1��Zär(Ǆ���Ղ��*�ฤf&H�㪓����)E�S�[-� ��!q�̜ϱB0	�Ir*�1���	^�LƊ�P�˹�8m�IH�����S��i���'?p $���5\�8�W2�7WPC*��JV�{��P��r��~/�ڤ��(��!+��l��*��MEqm�d*�5=wH�ON�KW�,�T��E�aZvhw;��ˆ�DQ�s�]�3�4�{Y���&��q�.V!����u�oό86>�ext����zJ�2�C�j��>