XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H���D��ʻ){(��4��iv�LX�6`�p�?�g�b�6�
�Ǿ 7\�D.9.i8�ӭ�q�V��3��7#h>�qR-"��L9�XehV��$#N�L�î_�=J��B���2��OE���7��\uu+c̪zVf��6"��B=m���n�Wk���!05�b�3o���8�VaX�3"����O�5�4��~Ϙ��w��n�m�C�	nE��!{x�	[��+�#����n*\�S��:v�ȋ ;G�7:2��Vny��m*�h'��?E��|��<ɷO�V���
d�'a?R�Srh!����E�$�?���^)�l�ָ��� R��2�\ך�NɽN'��m�!RO��#�J��;x�r���5��{ݓe�J˫��=Q޺�o����Jb�!�q�e�Oo,z}��Mh(\\·�u�	��u@,��� ��Xg�B8Z�oD�[	�Ջ5M�̞�a�ˤ]�c���c�~:�ڥ���G"�Q�Ŷ�i񟴏}�� ����uD�kJGi?�cH��{�"�����Z�O�C��SG<�� r�Jh+��C\��7�p�4,��Ћ�����������]����\ו~jG� P�t���@/�L0j�%�UЀQ�_2�P%[�6�����ۺB�m0�o���<���W�
<d�ӷ��
Ac�o��(�B)j1�Xc�vÿ@���"T�.�3����Pl)�in;�e�ˎB>�p��21��g꼗��,�4�ub����_�F�>�};�I��\�Fe��>XlxVHYEB     e07     680B��#EJ��3�S��\���A���cg#�7��F��6T3��)B����?J��4Zܘp5� X���[M��0�O��#��')�.-n2z�d���v��������.YC\����s�>���Δ��}��Bm��5���ĔN�n�h#�#�Y�wh�7�5�l�\��C����kR�*������3��(��?�0���4������EA��_���Gi	k��;[�:��o�X��n|<�WaV{
��ѧYI�z������qۊ�����k�w�TW��N��A����ƀ����B#"O�֑ ��x�^�0�f>ptm��E��JM����%���:�N��5�>���\�C��OH+�J�`��\N@�w���H���g��Ȇz?jL�}�6�4�JQ]:o �H���������3��t�NU݄�=c���U!�ԘJ���#}K_ SoR�MD�S��{�69�+������|@tp�j�Ԉ���"_��EC@�I���E=β��	Z5��z�����,P����=m�� ��>"�,U^ݰ0�59�Et�ŦMQ��g�����s��=7�D��E6��t7:�ϕ�d���xMq�?�֚�9���g+�	q��4�5df�������W�l�DR@�����f��tHa?����c��=�+�M��:��8��H��q�\���a��X�1}{���]W|�a�aמ�}�<�B�]�����ҹ3��,i��Zz�ك	���� A�*)5�ӪW[Z�Ě��Z�����`���ӑ��q�r��!����-�!,�wh�}�-�����������}SLJ��L#���e��(w"�t�^%K&�:@�<��՛��u@���;ɮ.�B�~>t�
� �c��G�'�gc	�pW}p��ao����\0#��L+�`-<� ��t7�F�y�����:=�P�O����ս!�y�Ώ�D�\�������tzx�5�tL��d�����%3�blP�A��Th���*(��������Ql�3�c�*�P���kG���J�B��(�_��4���8���Hʩ-x��(�;J�[���*z�`A-�{qB �g`���zᡦbD���o���v�y���ԅ�@�A��1� 69�H"��aJ�Thy���+��93���p�Ѥ>c}�n
֛G�n�uW�*-�:��rt!�AK�l�#  P3�:m@Q֨�&=�6�z7`�*��&��w�c�O��U�|���#�қ��,�q�r㰊M����7��+�$�y�e���s�w�n���m��9�#39%�*���P�nɂ�<l�I ��
�o�!!N��Cq�PFF,��)P)N����Մ��cDA�B;[�{n:4k%T�ڇ��cghҧ��EO��t� �x�>���z>\CF
�����s���FsC |Z���#����a�5n���+s��9�:�M�tv���P#[�F��w��V:��Z5b?��o��4�1�{�c<�y;ЎX����E|�[י߲w=T��I�:���?B�[�@��8��ω����Q �W��j�_�@Dj�*��ȼ=����; @f8���a��I�C޴
��߉�y�4����#7�w�o[�Ÿ��'{�}�f�����1N`��Ԇ���<�By�1*ЀЁ��ys0W@�%