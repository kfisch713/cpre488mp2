XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�Y߰%�ՠa�V����36l	\t��y�V��k��냤��P� ����5�����嚖x����|�M�吉�W��=a�"�VҠ>�֐�,#����YCC�ˁe�Pl�Ё�'��^I�D�9�Y�8�2V�Oz���sBC�|D0 ��ʣ��3�����N�p�cO�=}��u��уV��Dh�v?Z��!??�a(7Gh:Q�gL��yO9� �I�.�ʏ�C����m_G�Z5�u�A������~�u��Z��^a������b� �&"����sq649:�+5���RIH�KI�>��[+���'"O��e?���p�$H��|՞[W-me�k"o6㟜w�م)����;vr���:S�!S���?xd_Cf �ɀ��ƾ�ww�At]7��B3F����$������bkr�.�XZ�En�}�i1R���L��`ɞ��W�"�HD�b�j��Q73���͈n�����g�èF*��j�(���a�br���)�Y�IZf�su��Wd�j�����e{���E
Y*���Aw����ڢ+܊ �_ܹ}�f`����8~�(�E�r��ٻ ���\����	��`1�J ���k�o�E���'M����"�9���#�M'Fj�g,������g|��B��x��l�t
��禮��a�Φ���^J��/A���ؙ�ÌiΣ�1�X��z&`����b�u'4���:v��� �����eE"�)�-��plKE5Cx
��rO���V�XlxVHYEB    b087    2540���`�r�0�苺VǾ��F��0�*2L�'J���%�ɇpg�n�U��s��_ ֌4~d[��U,�$ƩfJ�Gl�m��:e�\.���ם�����S8�t�V�`�C � �02c|�PV��9�A�+>b����+����I�]���g�qk�<�2x>���(�d���E�[�0_ ���h�K�����W O��)S�@娨�!m\ab;�L����/d�0�o�y]Ф�	���8���}R�^���bt/,�"�~�$ۉZ8�lg��I�{6Tܮ.V�$����7qR�3�%Ĉ���Ψ$����[e��Ո�;��-5zV��M^��iݘ�&;aĪg�`��#�A} ��ҍ�� V�1����t+���,������v�� @M�s\O�ߩ������lm�L�¼~q.ݠ��M�*>�n��H�sZ�·Z��Ö�G���	]'/��^�79�|L�z�H�>ݵ��N��^�qT��av(l�X�KQ���BŊi*b�B��R��m�E�E�o�|]T]��բ�{��ٮ���K:��8�x�ɮ���kC��k��a�"���V�<�!���S��4��[e����S�U|~�C���y#��]�ʰ�M�E���9�;����-tӾh�4�0�*��#�9����6"�:�	����ׯ�b��=������dw�i}E��x�c�񸄧J�ec��&[���|T><Q���LW�L��`_�F�.��=�2�Ŧ��:����L�����n��Ȇ��|�y��A�VUU"��a�{��?R�a3d*��1�)��BƢ�aOU��H&)1�K+�Bk��7�h���z��vN^j��+���6�-M��-2l�՝��²�Oe�ӳ�0�C8�>�.��h+�����ⱉ/�^M�{'V�G8mc&�m�o��2���)b!�G|@�	9Ux#�k}��{�<9�qb��\n[U\�ty�J���Wq�C�I]�8MЅD�m���n�z�)&\{��U��%�v�����ˬ	��	����V	�0/Ҝ˗��|��CvC�u�w��P� �'��^̻'I�O����
��=c\�������D�)M�z���v�v/By�4&*y��9��p�
����CI�@������V���������.~t�"\o�+8�i��0 �()�����0�ˣ�"������<��2�h#A�V�P�P@�
x,>LVԸ��8b�G�"�E:-Cb8U�KPRΤF�,i�P���Nj��!	����F@�~���ɾ��n�����4.��48T���y/�Z�ò�n']�q�Fnǎ1S<��[FX�=��tJ�̀���`���-�"|��Y���({�����P�/GR�.��s���֙��@]���vPC"��<����`C��$w��$��~V<�=u�_�o��{�r}��k�O|u��gN���gv=�ȃ����Xʫq!�<^J�l��+ʼ���eI��cGr[�"�0n���r�]Mwı)��4�d3pP��n�]\Z�����a�_�1�`�M�?XG��ֲ�	�� ͐NVp��Z�����T���C�`�_�I��&g����*�	}V`�q������c��'6�M��D�&:=8�1��A"#b���^�#�\:�itr6�YLF=aVh���_i��1��vvz��<�a }��#�D��M�+V?
(
y��L?z���Q�YF,�@$�T
�h�d���R��:���б���h�E�=ѐ���Q.V�V� ���2Vk!~�i��ݎU�}#	{ �[D�]�k�%�ygm_z��9[_S)��p�:���L5�j�z��|���Lh��Ë͆�uD�p��($I�n"D����%��2��o��w��b����������$]B���w�]��xf��lXdC�HIw������*��7�[}>i�?n��r۶����u�"|�,p�(?Xו��]����kY���5$n�I�<]��E�\f>ˑ=%�������һ'�bC	@�0�\��'ɵ!��Gǉ�d��{�㇡7���;�����+�[��+oc)ۮj''�[XK��i-ȧ�����x8�'����T�T�eox�HAX;�I��?]|j��)V#uLo����j�Ϥ.k�r@��b�=�6}hi��#�"�B��u��i���oP5�0p���N`H+���=&��7kh��D�x2�	/T^ĀY�'�<H|��zt>�P���š�)����}���i�MC��3��[��jO�JQ���bمk-���>\P��E����u�"�0t�	όd��(.�+�Y�����pQ���|�ܼJ a���=_�n���!W�����̿i��t�l]d�*mQ�D��0]�v[5"��$3l� Xѓ�ޱ�6���܏� �g�_,�� ܷ�%����|�T.x�86��SJ0^�A˶��1+鲤��� .U���Y��.SY��Aꚵ�;
�M	L�^�J��j�`m����V����ǯ_��Q�T&�q��-2Nu�uz��Ն���w�����(�ʠL���p��)����G�G�P2'��Qj�bht�8D���:Y�^�]�ޢCn����˨�1��7'�C+���$y�޳�$J?F�%���پ�~|&7նF^4�=Z6��U8�c�Wn�}�������=��/���C^�	�z�? ���2��i#��~�z���� �~��/D���J��!;�A�z����Z\/���f8S{�~����O�?���LP��ݜ����BT:;Xլ�\<��$��fEk@���^�u�K:c��ɮ֒�/�K�_�����i0IM��}���R�A��ϪJa2�NT5��v�ND��W��a��"����m��Y G�[��\�������/��r�[�ڨ��ѥ�|S�P�򪦀�w�
��I��*A1�I<�+��Yp<.+��ƕQ6���?��T�<�h�2W�"����>�:�OQ�JR�� '��0�Dl1�0�4=Մ������R
�^����,U�� Cz�+VB��@P�#z�]���1���ц���Zb)�O��{��p���2��O�|0R���u�$����#fD����DQ̟�H76�4K��䏴T/|��ٌ&ӭv�]�e���Q2Pz%�X��;�i��f�E���*��o^+��B+�3��=�ѡ��P&������}���H�SJ1$���Ξ��@�f��=�����,Q"<��}A�MD4�6s�L&n*�k��N�-�/�����Y�m�}�QύH!��_}����m��Q��S�0�'����c���:�Y^q��1)���zp�R��Ǻ��#�(�aF�`�w�p��3��dQ/N��� q�[�R�d�9�f�0S�\ɰ���SG�ʫ���Fz����~J�߻j_�O$��= ���*A:���b���.G�Y~�z����oՙ�i���(ޠ"$�:.�S�n��\�⨁�JG�Q �J��)����.�����<	����`�0r�-|%6b1��D�fZ��(�ӄ�Mdi����j^�Xh�3�����5��f�*��vo�o�8�d�M*٧�(�;����,�������Z�SdȐ/^�VBv`��4ΆB��(8�' �UڎB/����W����E�� �a�5
����p��H��CHVw<�Q|��	4
	���l��y��_c��v+��ǺOY�/-�U�����`+L��X0L� G���gh@OQ4��Ǧ4<��cT�T�]�[ �%�{�VRʐ>"ȭ�Ѱ[5T����q��i��*O�.L%��ײ�C�=�	2���Y��5AQ�`�@�A<�	��L.L�{vd_-���X�v�����ְ�l�3�@�,Rk���Z-�}NmK"�&ޞ�7��MH�}� 9��ן-m�;��M">
��1�s"����&�ߑx�,P�Q��P��B�����I��W���p�#���&�j�Q�W]h�[�ÕO֮{�N��;�>��k�l�I�i{&�qL���q	QJ������������('ٲęL�]�z��{�LZR�A��t�q*
pt��Q69�]�hR�&�Xh��?��@�=}��dl�j}��F�t"i�����́[s7��p��2��D�!�8Y�啡E�	���∝�
�5�F]*�9���s��0x_S�:�J�{跺k`Qrg��6��Q|�2l�hMD;v�P՟oc�V¹�!��i�����#�£\���8+mi���lU�]#�{d�`/+Uzґ:n�q�[�>-Ǉ67޴�	�v3IzV���3 ���
�A�ϔ��)]P�$5�a���y��ݔ$fa"�>r9 wZb٤d����C#)ׄ	l+y�b媒��5��E��_T��lQ��X5��v/�?�U��i_����R_^eW{|��U��0Q�*�aOs$v�!�E������'��&I޴�f�ʔ����[N�=��'�k
�����~��,}u���~�<���w�>���������:#�H�XS�O�O�q]�2zO��2^��Z���κt' �C���/Z��}IN����aW�J[��l)7 �3���T{����Ɉ0t���]�m;X;��8|��-O��,��w �}ܪ�3	�b��:� ��7w#۶���'�/q���܌�1F� o҃uN��Y��5�@m<�L��]�U��'h��;����񷨰`�
�t_>A�����I,{�>5YH�2����<_CM�V�C�ؕ��Σ/���'1��P�'L/��,l�ţ��B�_��t��w_�&`%�s��@r�d���T<�7�NL��D�I��Rt������d�o��ۆ�߼�H[RQ@>6u�0��x��l@�!}W1���ɂA�B�g������F�G(V�B��7������DO��+h�R����X�`s���&�O����.��xǊ�q����;�˲91Uh�p����>��Ҥ�=�L���6��b��(�j��ȻA���k�����_X �6�e3��G��?sHP8����@�O��[:�;m�T��e.��{��m�����*�8/���TiJ=�޾������4o��7�d��,���e���3��I�|wJy�LHC�����墱%������.�5���R����_S4������L(��)^EH�� ���`�|��:��Z�t���*E��a
�Œj�J��	mα��Cc%��:eV��6]! �za����OsLSȏ��Q��h6�w]�2`���ΰ����B��`�82�VP�:~i��Z�/Ud�����G)��G��?[i:XI��K�d]�;��d!!�[vL</#��r�vQ��,�086�I�H����\ٗ���N�6�⋧Ȑ6��91��h}H���ڢ�>޵����K���� �%6�e�g�ړk��>���!Et ?3�N��.��^��O��;���#%�8�D�<�.G��*�%�~�~�=�z+�4�{�P0s��-�jpC��C�>�:5�v���\u�{\�uj_�	��8N)ˎ�u�I���<��I���s�u*,�U�;���I���E<����LC�ߒ"��(�0�ܪ�ԏ�6[8�BobAp/����)�Y��r� 0��ښ<���rN@A4;$�M�3R�2\���w�����1��Yؤ��8pX��$]g'�>�AB�S�=-ŧ�M�Vs��>ިt�=���)��Ak��k*c��g�S@��M��ݢ<����7,~�p���
�#4�=XЊ{����6T�:8\Nf͋~B�ms{����m�{H�ӂ��9rA�����3���m8�L=���w-����ӯN�s��a$OLM�5X��M�.��-P�r-ۨ�yK�BݛW�E�2�O񄾹z2���{���ɛ�s�x�������1k�e�p��gh����G��2w���q0�tp�����6�⣒���U)E�5��9bP�LY��e��,l�<L�VJ?h��~WG�M�a[[� 8��0w'�L�e���!DZ`����p�7|��&j�F�O��� 9s�C�-�1�Q] |���X�W]C�]n&��0�#�
g<pGԿ[)�y�J�����PH���[�,�ǜ5�t�U���cd�r�X�r�B�͸���n[ ��H"g�Q8�
1���-x��T�����k΁F) �L<{n���(�:1(M��=_� 3���i��'��#��(�� ���uo'I�uJ�I�8а��tR
����#���c�]r9Lݛ��sj�Â���+n�'C�:��>6�!Wt�v�;]+�of��B0I�D;����h/"���T��:�)(=��
�o�K�s��W�6�'�D5k��[x)y|�0�؋�T���i�i��O��'�hvH\SA�K�l	[�{���Зe��.SS,"�
Gc��J4}�����3���������B���rpD��"w4�۩Bi�]�I�%�"�tk�+iU����m��)Z~n"-��t����.�s��<��a
nuT= y���f��ưf��f"���k����3R��VZ���VÞ-��6���j_8jL6�Ю��s�*hψm��h`�5��LM0�=׭�**���]�o/�=~*�.ݮtiwV.�y�n��%Ҷ����|1�����lEDZK���eׄ�
{��0<�_��=�5�6�(>��IЌ(W�sy�Pet��!I��.���L�'�,����e>BYK�j�=��IWS���!��o=���f���`��Y!����|z�0�=%�$w~Z+�fV8���g���Ә&P����x�jsI�U�0]y.,ng��iI�7i���T5R!�\���6:��R�̰��r�_iU�]�~>��%����������y�u`��qb���5��0��
?�2�/���a:�:�uVQ�b�����K�L���F�C$H����W��(�f�yk����I#���Y�������䓖]�8r>u+�b
�t����l��,�����?��ʜ��b�0�("HDnfhRk�"�M�lWe��o��'%�KC�[�/��˴���s
�A��Ȓ���2b&b� r���<K�Gb�2�z����G�I����I+��G=�F��d_A]dd���:���@W<�1U�dS
�.���8Y�g�y�?��@�⸃�!����i���4;�K�uq�SO��t�x��6����������!�f|Q�R� �z3L�?v
\���~B@�Ⱒ�_�����R5�]��Cg�������,���g�.5� |��7�lء��^'@6�����0�C;�zMiE������XI)�D]�`�} ��H�@��^.�NY>��"�p�n#I�U���=G�)��!qj�ye��ug𳃲�QE�'9Y���Y�nxl'.�?���g�H�9
�$xV�~���l5��P�im��9�҈���[w�)S�e*Z�b��{�V:'�]��_����`�T����ʖP�1g����!�,c�
�Yԗ_f�z�&�W��@���d�ket%7F?۩��C���uc���'�*m/�@�d��;.c	3Cj�WsS�6i��#?���	��l���kP�f��
\���ά�B��;쌇O��!�������f��G�� 3�h��VVM�O|�!kb�����E�D8��b8�Vqn�[y�<��}��L-��+�Kv�`)��'Y%��B�g��iw�c�穚��=H���/:�����0����xV!�\?+��g� �mXA��tX\PK�5�-��ǫ?Y9�d�u_�B��r�7�IPB��q�Q��?53���X����$FcӀ75�W���}��\��_�s6𲜨�@�Oy�9L�Ix�� �O���'Xk�)G�%d�"v*��2��Y7؉E~���HuD���1jeH����`��UE��T��ʁ����e%��ҿ������F���\�<���_�gcw�Zb��Vr$�֜3�'�e��N�!�����lC]���=������]�z]L��+�Oz��cT�A�B�*
��Ȱ�{T09<�g�>L�LM���?!���Ꞩp�Ҵvs���V����뚖�5��z�T���k� ������P�P#}{?k���� H���11��beW�m��:�3a�sM]�0����o��6/����a��3G
��6�`�b9��a��� S=�z;��.S�T�>��B�����ٖ�\�`�*��J�g���|��� �/A�*p�qt�`�&K��]��e�a�YC��ZnА�iɨ��J���ǫ(�rh$E&-9��ۚ!Cz �5�ۀ��ͩl���G�5ڦ�m;:ҹ�ZN�94R$��Dw}��j�7��g�Pm�!ġ��*A��IQ?xrX����ի�:�R�Z|R��pP��R(�N�X�ݢ�,��9x����|�4Tk�<<���t��2|k9c����C5&�a{�uC+��F[%�+Q+��V��b�$!뙗��f��my��6���MQ+i���d1{ts�9^���z2��ڸ=��<b�Vօݝ�"��,�_d=�j��nꄠ�g˿ޚ����`�*��|g��d���Ӑ�I�7#�C��s��k�#����X������=!&�|2�a�9��@��8�4eJ�eC߂����$�5A8���}�̥�8����MT��3�lm�""�Cm��(��Y��g'��"<_N;�@�*�*�#8�&^���d�����Ns}N�O�j�Nc���3�'k��\�)評�G�˅NK0P���q�[�H�\`���g�[�:�"L�t�Q����i"N=��-6ښ��@i�͘�р<���e!�`�䫟K�Ȝ:�V,���������&>We�Yy�p��.������L�"]���z�����b����\.o��O?��B��?S�l��v�Ⱥ-���:���cQ{a�=��7D�Qn<9�.�{rHI	���4�-K6oY�+/r-!����=O�-U�,�7ƧbZ -�X¢~ ��k�3O%-�����R�D�ܺfxp���{'��6jttSЦ����0xM��J�	K�^5~��$)-�g�vp����Qk7e��$�=�1d���]��y<ރKg'��8�LɩŸP5�>	QJ����s�\t���U�OYjͱ��Y,u8 �9VG�K�([=aGC�M���j�{�Hv���j�4��J��M�|*�Ӟ/9�Dv��F�ޕ���$/o ߟ|���2c�^�`��7��+��%��r6�Jh�.9�E���z��9x�����^]2���aʙ����r���ݜ�e���wӌ\N?2�v�ǌ���}�[*��"�ψ���d�e�>4�