XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��nsh�^�N��?�^�X�K�Mo�鹤�I
L��?�f�=+<5��2F�˟�"'hT`ӟ��I�9�O{�80	�:�����'ٶ?��D�c"�J;U���(��2F$�p���W����NCNY�]_x�3�����b�iE�*�����"�h�0�V�M`�~"�Ř��jv�?m}��؛�p��p����r�4�x(���"�׽7cF���ȓ�_]��'�iLͲas�]3H$� o�z��V@��ZKP��I��x�����[ߪ�[ժF+����n�� ,�~,��5�J���f���?�wx|6�,�0�ڮyq�b����󜊍�t��d�EO�C����W0����G�Ч������dF #��������T��Ӫ�ni���1����M�*4�~�B9zP[P-5PW,Na���vl+&�{�z L�[cy�{A���G�`yU{�hwӋ���Y����7��솾�+(/ �QK�6���i��%��:�y*�'�0�3;�
� M�~&5.����D�FZw�F�*���'�@ͥl$R���ilea��t�'a1&|I��C�l�D�W�S^���>���|�-�#$\��%�ᤣ��s=��[Q�:i�0Rv:��\�࣓7�O ͯ`ߓ�U�4ftI�>�cM�� ��Qx���)D�� ��,������]	{Ρ�wS��5��0�ܷ��/յ�t.�+O�P��D����z�^-T�}qϒ��B��ݿ�'yn���qVJT�����ڥF���XlxVHYEB    15bf     890�;_�kag18��)~78�A-�?�Ys؇$2�@}i2���"d�EQh�����q2����6����DS2�n�2��lꤢ�""E�)���4� �A�B0��24�oG��
�(���P�$.�Z�;��D�0g��.lK������Z��A�w���ډV��z���ν�RU�5I~Py�1���/R�@��#�R�Zt�j����|�Q�9=:w����6]߃���s�,��'SF=������������rX���?��
(��Y�l���\�Lt�(�d1��H��>V�#���%��B*9��F>C��xw(v�{�{Ƕ�G�$��{��f#�d�,�# �&�q���l1<�N�> �j�b4�
5��8ň���sG��t��9F_�s���c�m{�J�葉J��s�(���?��[L{0��T�c���^�ݓFA/Դ��5��0� !�з�@�b�~�	P�6pBz����n<�{Tl��a�rq���aF$�A-!«%��<��'ē_
H/0���z`������	��X&��t��+���	�����o���J�*���Y�Y:��\��#�q|?H��Wv���:�!�PLΌ�����zĘU�^����2�6#e��@��>��?��:�̜*����w`d�T��qfe�&�֡��'�J�h5���39�L�p�׺(;2�LZ��{0og2�0�=i�@�� �E[R��D���h���;���� .��ʩ�`e�O��f���N[t0��u�X�	��؇�7��ͩ�b��O�n�� ��Y���T����5�J�����[�KO�Yhs>�3\�������[�f�^��r��4B�`���ŝ���@Vh~��Q��:s֘VW�8{]���Տ��h�jgR����'���� "��l�b6�)�ܙe���		��0��NI�+Hz@ؓŵA�m瑣Ҋc2��؇1Xp����u��������{) ��u��ZL9i�m�n�X���$g����W��k�R�e�I%��Fq�8����=��J.o/�Tn2�YT6U���1�-��;Ua�0�!�}ki&�����M�x���U���{S���-�P�HPw��g���َ@'����W�E!��O��o�m��i����2��KKೃ��3k�N���$�@�̍1�׮ؼJ�LM�nϴ��Y�d�|���Er[8������5?3���N��� p0=T���K#߿q^�I
Q����=�B�ϴ'��!X�*���' ��5M��פ�A`�(v��%&�v��B2l�6��@x\�w��j�<����32�M�t���V7��6p&\;E�K���r�O��69Cj��U�j���ylP� `LASp|��xlf�33r�ΪE��r
������OL�~b�^�T#;s֗�EuA����}�&e���<�|��d]�(��nO	�8�Ǹh�|���p`��dQ�=��P�)���Ѷ�G�x��T�=[Z;V1%���qKJg%�����"^C�ޮl�f̣@��o��pZ��lF�4̠sQ�-���wb������m�2�����j��ё�2�eP�1�����Lm�"�$P=��=ä��ON�Ǉ.�4cR��$x��a��w��8L���DV�hé$DP�=��w�:�$�X$�F���X�s^���5�C�I�5h�9�x��P�Z�g(�@c��˹���/�=��Q4o���}0��i�s��MJ|8��/��ɨYڞ\�'�硖�[�yq2�M%΃ͺ�W�=Fnl\5��"W�AL�t��Po^�+`��P���F�m���	��������s�e��e��!(6}0�Y^�'c@�)��+�`�0IN՜3�n%x[l�K@�+r��:��:�0$}�#���[CSy�X��Y�Y�L���_�Q�@�`�1x�V��QÍ�9�s�r�)�#�����N�5:��*RV�ȮS?JGv��F��+1Q�Μ�L��
���I���,:;��9�ն�̮�=����t�1���D3znJW�j̀��z_)A�> �sI����{�ٻ�}�X�;�C)��>ЁD�yZ�'��wӫ�u^�����xWdLce�2�
��(=ݧ|��`C"�!�����i����\ �3 ~A|�?�
��?0y���e�