XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����͆%�lnN�p-�H��k�&㪀&OxD��ʓi��'łI�4k>�!��7��IG����F�QS��px�8�6��k� "8�#<�Pܳ�q����3�_o�t�F�"nw: ��#G'E�qB����9��giJ��
 �)<+�Š��J�D�Ǐ]��&�>	��0�b��ʂ:a�3C�c�Vܣ�ٱ�4�iic`��?dIT�ޥ���w{:)J����V�kR�}�9�ou�AS�����OG�g&y����^^ek6�4�w \'��t�ϟ��e���eK��~M.�S�L�T}@��n1ۯi�,|0v�A�w<ϩ� @��O��ߜ������5� Y�E�3zRD�q a�)��dr�xE�7.���E��ɀQ�nc;�3H�^KBS�a��b�pZ,�_W�<�`�V�-S](�3{~̢�:%�Y>����~p�޸;�������l	k�+G�R��=q^Pt5Y���2?�]���Z�E�	�s� 3� �� 8�굃7�H�J�� ��y�BJ��e�L�A2�=��JƩ���և5����Ҹ����t�^�_\��6�J�ix�Z��t��?�l�ǒ��Ѽ�� ���8�3���/'�CS�
=<FЈ#��$�A����:�ֺ�<�2��'�����A�dhT�j�=Pz��7�HI��VkV_�>���K��`xi��vHpAo�+�t��L��nCs.�4a�0��
0��K��J��ةg�0ev��qq)�fXlxVHYEB    3b09     f80i.ڗX�M��X ��דhK`�4��ݛR������(�iM���v��;[�de���&D�?�������N�M�3��F\A����?��n\^ȫF��ϡ愃n��7�k�6)|}rJ͸6deB��7d��"�?(1�ɞ#�s�x"��QcK:1gcڭ�n��K=���&O�����;r᮪ݨ�c��7�7��0<���H�w�uQ�w�8���*Y�S�0ؤ}6�M΄o�3�i�@1Zޥ%�a�g0�c�0]g^+.���22�7Q==�q���Ki�X��7)�n�K�9��"��� v��I�w�,��7==�C�w@����RXpl
#{xX��v����:Y?#D���HV#� �Ч���t�G(_5���75J�P�\�+��w��E�D9ɲ��#�_ա���X��OCL�o\�-���!�=��l�_����ۗ��I5߈S:F���OH��NU��� ��� G�+��a�au3�f㡚��g8L헊���n�m�(8�	�[�����dXm��T
{[����,��n^�լ����y�(�,5��WhZ���~��@BNgJm6}��	�}x��όE���/�Y��]ݏ�%?ϽZK���+zW�#|�]��4��q�����
fS��x���ȸ�"0��$A!2�]\7b
���}��e�"Ъ�B�7٫���c_Q����;�B������PN|7����p}�	ǡ��;R��rMk�(#�J<�\}�_��p�4�7���6?�
�2k�Ǉ4��Ca(]�W^Ax������(�M
���'
jѢ�Z�S����1DX���9vg}K���mf�$Q1�n�.�袰'J����C��hٟ�Fc}��f�2�A#^�޽)R>�*�.8̍���p��!S�0E9~kb����HyW�T*��y�m|\�ٻ�o�C�(�f�����Q�C��w���~���6M�{���'���{��'m���Ou�\:��@��l�Y;w�
1	���
4X��5B��
�=]�����g|a������5%��� t���^��בS��N߆�pa�z�8�����E�[ bw?S��.�����}��E��$]�ߖC�/|S)����;$N�	�T>s|���}U��C8k谅�+h����`Ud���\�n���צJ2
M�h�ؖE-yY�;�)��&�^���Ѡl��ŐN�G�}Ո�f�~���'�D�P�)7mHZ��BrPr�#�ge�$l�
n�a��!"�f�S�;p�ѫO�,2��&�,k�n��KvI�?wyU����4��[�\�/�wI���;;�\�:VZԴ��3��' �±��<�R�w)jb��x5LwK�=3�S鏰zs���� q?�#��/�1��dp�m&`*2�ֵF������WaҠ��_��8�G�v�d;��m},��暉(�$>`��nȺ����c�x�[�BF��Х6��o E���u|�d�:n�{%��C�~J�"Q���JF���I�YR�Gn�ͦrA�ɋ�Y��+uGb�R� t�����������]��0���co�y��Z�F����%�qCy �R���7��b\洃�n��O�2N�tt��JN�t�Ʊ�iF�DIT)��|��qQ��Ц�}��;�e ���4p�/@�Q�����9<j���l�(��͜�;˕��:��y��q*��ޔ��a+���p[ �I���DW'��Z��]�.�R�|�%�������=H�NI3���3Ē��G��0h}8�f���'ᬾh���Wq�tMpV9���ϡ�e���]��s� nL6P<^1:�xm������t��r貫ԃ�$)����zT�O��zh&RHKh$�/a��4�Q��S�5�ԭ����E�s���N[w�(�<�ՙ־=�i>��BdP�ߖ�d��I6�����8=��|vC)�H�$�'��'��k�@�uL��d�ŖY>��q�x!�B�y�*��Ǭz�݌S̕X�<���JH3\� �Հ@K��UCc�l��%>OR�ʬ轍ǣ>c.����|�V����P����{�����(ͅ��ԣ?< ~B��WN+��׿
U5i)#�8b� ��Q���+d��8�vD��lݗ��h��Q���E�U�D��ɤY�%��[�RjhS���}q�
9�V4Չ���D~��ց�\���S�>���F��ȏ�u����5䗇ؚ�����lJUL�ڎ%B3"_2z�hQ�����P�Ӓ�a�eCy)�]f��vhk������y���u��O:�x��M2��4Rt�1ˮ(רOxF'd�2=��KT�Hp�+����;G��g�����;�����^�b�I~�Q^6���$"iK`w
�x�UB)��w��V�2E�lZ��6BJ����D�>M�:��ý��oh?7��bf��A�,��oޭ�����%c�1�~?�@��|�c���^�ֈS�����ɜ�mVtf$1nAn�§�v3���� '���ص�!jr���k�-Y�P��H���^^�����'�1!���m�u*7�"f��$����N�; �>D�8*��L��LYt���J%���"Zf�Sr�l��r�Ü�؏�\��"aܙ�ߍ��)���H�c�Z�����
��[�_nMS�9ꁶH�2�_Ӵѵ.�7�n!�V��k�Gm�r������av��ؐ����UtZJ�8��S
K���݇�EUŨW=ɔO�l#�����v|KG1�j �7���ȭO"'��s7��ޢ;m����@�`oh����{V6^A�%}�%|����Т�'-��{�1Ӆ*�$}���U(�=j@��ԅ����Oc$QUEk2�x�\OD�)�ݵ45|�������V��(�U�Qj(d����y��kPOBʁ�-xd��o��4(��]ua\�9��VExw#[wЀ{�S�.��4Y���e���Y��yZ��'�Y|���=�)tj6��=T����x�/4���{��K۳]��=�@�ϱ����n�,��
}ʛҝ[��
�ϕ�Ss��a� a����A�m���(�ED���wK�T\�<��C����HѶה��AB�[����s���LY69�?z�P8�=V҈Z8:%�l�r!�=���#����Cg�)�R,]�d��p��u�9>��I%(��y��X��6��KJ�:�%������]������;rZq�@'���V��	Z�bXe��������?�#��pޖ#�y-~8��jF�WR�}�`v�ԉp��qk��=z�
�C=\.l��Q6�d5<=�P��r�S��=�Ճ�BiKl�/8"�?�	���1U�5�EA�ՒK�nKM�$D�=�[|��Ƴ�A�~K����W��+#�P�2�����/=�cC�`ȃ��0�[�@��M�8�a���:JI���G��U�Q�4��qU����x�t_|_����Z�u��]���z�a��&�*em�W�#�Y ��tNFI�����.�<���J�-m�(���lM�������\�9�t��45<����TP�����O�ڃ���ҵ���(�to�{��h�!�y\�y�7��#jP��g���d��j?7�S6�������(���18��B���{z:���~X�rt:�I9;������ĥbu=µ:3���~����*��[Q�ۺnm�v���5�:\H�jiCj�_7s������š��x�#��L'E���p]����Y9�g��������N>�/{�ZX�de�I�7d����I�Id#����ǭ��D{��F�����KX�@�dɤ`i��K�#=�Fۃ7>�X������t��D��������Z0�5��ӸJx�S�j�<�ڣ�u����b̓$�H�ݬ�;���eL���d=�&