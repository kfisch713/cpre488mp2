XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&�Zl�O��R<�j�ޟ2y ˆ�rj�A�+�w�Jr�|���^.����?�-(c���\d�p�-��@oP癪�\l�� ��'�{��&o%�Z��5M�\�P���)\�B~�x��5��jJ�VC�gح2_
"}/��P�i�ܶ�Q�UX�k��>y��S3T�	{��� ��L�B[�Q٬��Fi&��7_������sN|[a�$�ڕ���Έ(���F����� � �Ȯ��(��F)��s7�պ{bߑ1u���8�m��un�LCW��(�6P�5�V��Gך�E��e�`��o� k����\��.��xG������[� :衵�m����^iѥ�(!��`2��c4/�=�.��nʫ�ީ�5�OU���'�Z�3mXݡ��G��
��5�m�
~@��?G�<�ث��vᒿ�g&�go���A��Dܣ��M�Z���(ad��t��ܰF�'���Ψ@��H���rx�����˃���i�g��V`	��-Cr�X���~E�&?��c��y¢����2�ur[��-H��i�����l�������>
����ߌoG6� ��~��`�oU���K^�mD�Śx�����&v2Q��R!t�G���r�Y��Xg�����gS<�o%E0������Ť6:͏��+�6N*��Z�՜F) tʣ�7�ȫޑn�a0����1{d�%
'�D�b�=� ߩ1����2���g�De�F;f���Ed����XlxVHYEB    4b9c    1300<��lH/�X�$��f���߸�c(��2�iԟw��\�s���٭���*�4b#�t�v���䟻����'7�����TБAʒ�Eš�NQ�ԫ�q��{^ݩ+gw�K��<�#�4���jN_��] _F0"9��f�{uKB/ϋ(*V��7e%��P''Q�d�(Թ��`���@)��"�p��B�� �ND���n���&u9�([5���YZ�q�GK���UA���T@H:�T���A�����}&#���+��[�d.�F��¥���$¹�Z����u=1~�o��(�%3G��iD�$�����jMM]��E#6u�����$���@��.9��){��F^�s6�gǒ����!�LmvW�
����^ ��[R�z�����k�s��9jy�`�[�a�~�~� �����*�������z1x�AiwS%D<�����F����5���|9ȕ�M ��3Pp78��q��
�OV�&����4�z5T�Ci]��<� _��M�Qn���K.��>
�m��W�6��Oo�9���������ڈ���og�E����8�;h{$;��{�?�qv���a1�`��6s�U f�΂5A<�̈́��5p@#�5��<�����X!��1Ag����Z3����ԑ�#4�E��1�i\	�X^h���a"�K���WV��7�e�u���Z�q�:�|��u ��P�S��x�Ę��Y!y�B��]/ݖ�� �cPs���P��_�m5���v|�M���=R����bua�YE�nO�����[7A�>�?��`�:e�����dt��0&� 	U(�7����0wh�-5<|�<�\2���^{8�Mقc ��kJcH`�c4u�j�\Յ��I-�o��^}�n��	��z�J���4�\3�e쵁Ct��x��0A��t	g�Uө�:ƒ-N����$�-
#�B�����'���Q�ڭ����RT��d"�:*;���ꁛ�Ñ
2G��=�`�łG$b��$�j���z�Bm��O�}�Fi�vft.���B��[QE	��qxm�W�@�BK�4�J.����L��V�[΄k
�9]�c��d\;�4^B՛P���$}.��ԏ�p\���J�y!�%�Y�İ���L?D�ߩ��I�|��Qe����ޭ!#�Ճ�C�FцS+P�֢��3��_�Ķ��ϭc/_(��ὓM�i�VS�U�t��{�է���'��'F�B�������6�_�X���?4/mD4Ze�IKx=a�z@4[ؑQ|����cZع�{��r��~�C��l#��E�]w�G��X�xL s� 6[6������}\����t�A��^9�*P(����e5kp���;�E��x4�ٔ\v7���wδ'98l?e�Uw!�?�|������`�jp��4����B"?�aR+�c���^�YĂ��W�R�W����,���������Z�f;F�S�Z7�\@�!R����n0?�-��^����j�:N]�Jt�ɱ:��M��]�+�+x�e���3c���˦(�� ��\E�)�1����L3;9̴��W�W�������xֈ"���>�5Ӷ�n�ׄ�MW��ģ�%2d�fdFlR?�M5�/T
L�jf��'dmj�]���E*�]{��"m���r︳�<9{=�����ї�e���i7�SKpy	jᱚZ޾�i��z��t�)����{9��PF�2��x6�`���aҨ۬�-���Iko1I�7�ك
�"�p2�Rh{nl�������W����L�l��Y�o�M�ϳ�5���s�sE�}E��گ+m����b����D�bŦE���+��#ۚ{Q`��#P�ÒR@�q�fS����BCl�ӆ��`Y�G��P,�U)3P�����!<���K��9 �%y��c^��N|Ѓ��	V{e`J�X�*_��n���+�&��u]إ�X	;�j"E"]tQH�,U*Y�j��+����s�G�#����^k�?A��}0r���9�>�s�f%����
�L0Q-_q����,i�}�IU��ܐ��!/��s͚�S1��g{e���kL���S���8� Gg���K�L�Cֺ���Zgm�1��Y�"�x�1��(g�_���L2��a�������P�ӷ<��KS~Cv?d�������(I�o�eB;�i:�czj�j``@{� 	�
�Ѣ	�3ZhA�� �9�����������Ɛpҍ�AH��Fl?�ZN1�����x.
?VP?� ��|_3�W��������hy�U��EH7�vK��V�k���9D�7%��;-�/�w�A�ծ�y��C2�m�+����/�j���/�,d�L�5j�v[X���c����],Vk�<矣��M���QGR�ln"��Z���|y!�����I��˯4e|b{��ϩ ?�m)l����{�w��ЗVo���XO�����ǧ��n�I��%�]0b�ը�^ku쯎G2�7(�� 7yY[m.�rް5��	2�k�~���A���5X�{��S���+]��S�'ɇv���:��C�!KQ%����|1o�A����@�"YKz~,#o�&veȂr*3�[�W�mC������5���#�%�����u��_��E�Ln�\Y���&QX �eO�uG�]P����(To�6���O��4Ѽ���yQdJ�b�k�gw.�O�#7�<C�n�E�G�
ܟ�� ?��_>򩁈esF�!YXj��_��.����a���ȅ����S1���I5,x�|��Nx��D_��H�xӤ>{�Ƥo�7�2���o��-E{��"�ӆbՋ��T�����Yf��^��z��U���2��G���.������,
J��Dp.`���F�1�4����<���;����|�l6���44��T��RKgCl(/[3LyJiV�Z��8��?�'Yu7+N>��)��p��2@�0	��ǷM�O��!o �g��c��^$��<���wAG�bo[*Zau��S����������<,��?������}_�u?� i�]�G��*�����m��g��{���]ى���V��𠣕�+��V	}�Oz�O�� ���e���~��?��(-4!c?Z�a6�H��pz[�1�(�K��f��r�-��k7,��#��In�I��+�.��J�l������@B��TT���W��ǆ��w-`�-�/`>�ZRw� Nʦ����	�2s�0��GS������RY�;�_3�y��fTZ�*�L�й�90�j	�����tͩ~�pˈ��1_#{�k����w������c`���ޡ#�u�1�2�q@��U�_|�֜��Թ��W1L����A[�5.��<����8�Z��&��S-�$���̃��_���@�z�n.�kUGfW#�O�������z����4��I>ށ�||i�g�������zn�lâ���<'��-:9�TF#R�1��E�f=&����|w==@��q��j�
K��/�,tXB�OÙ3���dw�9K�͍o��Mp�q���)姻�Pǜ�j��ߡw6�p��І1u�cPg@�M'���`���"Y�Y�����Gz���ߐ�\�*tlU�Ho9>����vr�"4c�6~���E���&}lW��5���n��+��F/{��;`SN��5��ڴjnF6'O�#"��v�䙥�"`��2)@�q�t0�^�A��T�Ț��֦��DԘr���7�*�97R)��e}oOC�@�1������s��^,PS���0_��~g瘶��B���`3"�Ĕ��嗨h�����!0������Z�E��hukL��iE���9���O�8�j���aw���(Y����}���-�BzHs^|6�V�ptK�<���z9U��V����'��e�"N��_%�H������#u�f" ��F�jLO�ٌy�����`��"��)� ��.�uA��r�bs��FL�VE�H����ELԈ��ݱ�*�e{P�vg���95����!���j�OQ�`ڒ����w�y���	��)R?o�$�Ic4�������bm�G��.�yS��P:
iHNam�S�38Y��;%0�8�^J^���0�OEY������1��<5�>��Dn�mP��l��kh��N��� V^2'�T(�C�����8�G7�*��
���� �ܡ����FT��z���H�Rd����z��߆-�8��Ե��xT�"�Օ�%;2�8�zx����
��VDu�yG�}^�w�7�����<W ��\�$Y;�ɽ3蠓��FY�83�h�#+	�ˏ/E�+�Q�*t.�+�H���r/~FB�5�ta2ߢ`dznQ���=��d9ةkp�(�9���E����� ���b=���=C3}U�u)����-*����~�7�)�Rf��5	Ұ�X��]�������v�G`�f1�iA2� s�7��Sٰ� �DR~�sܩY�a
������LE�	_!��{ݛ��7�'��(��ܣ/�3�H�v�[Z��V��Q�+MiS3�ϓ��}�[�W-j?O5�O�9dC|�s�fG5Grh܎ z&�7��hY���tIwbW���n:ϛ5
ߖ*�F=��:ǔr�'�C��4���?�9���?ϐ���}�(�ok7���n�A[&���_�D]"o�*W?���n�(
�f��/~�}H�@>��jT����&4f֡\pq9<���������X9th�y_���"^C�I)B7�b�v�}W�m�R�S�����_;�%�s���@Z|���TviyB�f��!s|�