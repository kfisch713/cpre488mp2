XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<K�e������`A.y�r��(P�r�3%^qAyk�v�������圆0�|;k�������X���|u^��o�Jh��8p��ٸ\,L-�{t�*���0��Q����E�3��x� ���T�a��=\�����|6�c2���m����]SEll�AWN��m}��RkeKk�а�k��ׁ�SB,B���%�ep�-5��'�RF
Oh�#3�r�<p�7�Bx��8<t&��q5��AE�0�H��,O$�Q�b(�4���2o�xf��NI,\Yt䆅�-FW|��_��@;�֤U����Ë:���Q�M�Gdz��Ѡ�=�C��ǼlHi'�N�G�\ ��׏�2����d^!��b��R[������E������kq>� kp��U������6�7��JK�3~x��3*���In±!�����^��x�ݹ�.^m�B5��:P��]iǬe&��aTK�zZ��Io�N�D=�@z�cn�a1�1�4KT��ư��6���x&pҶ��t~thR�r>�^y�c����igZ��Z���r�)=Pԑ����S^']�ށ�E���	RD��lU"��1� a��2>|��	���~%v��X����c{q!�!��K;����2\us�I.c׈\D��ex�e��w���-���q�
XBc$�������w��,��	0�).���h�	��aM���0!�Eg>_c8	�$�z�G�w��I���g8?�u�����EwMO�0Hl��#XlxVHYEB    1e3a     a20�G�GL��{ vuo>��M�5���Mvߎ�hHƵ#��aZ�Q����Dvy�Ǳ��;ڧ���5ϢV ��v���+���ω�m��E��8bx�g'�A�o9�%ҙ��#�\b��2C�uO�v�h2PȖ�R�#Ǖ'W�*�f�b�#?��D�;�Ҳ���Y�y���Z�"p#g�IG<㍹e�������v|���"THN��U�����H4���7PUȼ���͇r��:�r���Cy�=�h�:ҵ�V�81#n>�<C��
X�Z�(.���ݛ�&F})B<-	}�C� ���12�SLy�jQ�WZ��i@���*#�Ub g��:4]�*|kȅ����28j�݋�gz��$�q��0�<�չ����T�5���:s|�GW_~�s]>EW��8x��{�l�C�ce�!�j�_����CPʮ�U\ަ�]|L�@2
�N�A}�OW����+��C�������ʯLR`��Xy� �p�h��wx�Br7�/UW>�[i?b<�	چ�\�!���q��}}�����/��߭Q��y<�=8fP����<$oH���D�� �owgCX�K��?:�
�.�G:.���;#��F�����G$kJ4��s!��=A�P9Vh.<2f�S3�ꜹ�Ɉ�Q�I;U@�Ƣ�p����c0M��o��Il#���D<)ͫ�C�� �kY��[���%�z��z�ghr�Ri#�����Y)Tç��s؏��HG)���߷2�F��Ԩ{�g�88�>ku)�/[�A��{п�(������t�����x&iO�i��U_L-�32�5Tf�rjAB�8�|j��ۿi9J�U��+@g�);z=G�
�z�qg�^�.��o�����N.Rc6�B2�):�D~���X������!����<���J�{�(Ԙ5�4Kx�<��C��c�� �q�J����Fj��CPg5H��B�5G����R�%?����H��ֱ�*��5)���3��R4�[l�zg����jb������oan'�a�K��Zk�f���+[�۽7������j�=�Y�r庹$<�q�����iE��V�#�B6Y�;��3���;R�D:	B������Z;�t3���������Μ��8����<L�H%*0 ��6uڤ��0R/Ff������?5���ׯΎ���!3��#�}x�{�zj��ߞG'r�i�TUP��hCܩn|��HaY�Y��C��F�E.��a�L�N�l��	���~׸��v5�ZEKƠ�W�F��_.��ӴSUN)��7�����6�.������i�~�9+�����-�_,�=��Ǵ۬�|���v�*y�O�Ü�Ik�ۀ7+�al��V��6�ǜ�I&hs���Yھd+b�!uI/��_�I�[,%b�j�����_G��ͩ�������Ħ�ĹZoкS6	�k�5�.j�J��k젪6��yi�l-u*�f,r���H�3���WV�|{�e�a`g9T��6P��N��;��GO�Hy���sp�|�A$��۷��M)���Ҋ�����+��m��CB^˗����@k�y�Q�7�w嬺i%Q^�7
�:�2[��?�T��7��M I
K ^���/�l�R)��?@��x�,ޅ93��隸�^������w�Ū��;�5�d�e ����ԩS�����E���ܠ� H�˛�Fi��K��YK��1Q��	�ȯ����Y�z�e�4�t�hR��� ���rX3��3�3/��t�2	�/e5d�j��C�ݿU�K�>pE�����?�a1�>���UE�F��b<�pG�:ʽ��H�1b�PjTf�7���-De�)Y��J\���i����t!Q8���+���T|�GxL��� hh	���yJ�.u͐:�� G�aw ���{e��ә�(Ux��BJU�������M0Q��kI�A�b?"N�u��j?@�4Z�-!m�H0���~`�_���q�]D`΅���N�j�x�E'R-��#<�]�5�&O���^�[[g��%˕�� vR�31&R�9�A���s�K��h�vw�h�׸~�O�sd�@�yQ���l�]��M�ó�X��U�b�L胭Q����� 5���S,�(]sE�ゟM����Գ'�x��M(��1Z�F�]fW��g�c��Q,]:�	�I�C�23���L6չ
��kz6�!V�緶�wV�{Ʒ��ͽ)��&\ʛIY� �Oh�D�B־-����Q�l}y�q�)��$���Y7W0����ŉU�NuQ��J�ך3�_DNt-�"�+}�I֮�7�����2T�6`�p>=Q����AmK[�+���r����B$b^�8H�#������X��B��xZ�x<�!N��S�m|�H�R�S��ͨ�1q�r{���#�'�.C7���PQ*��_��*<	ם�Y����r#"b$�
`݇z��u"�l���O�^i(� %ݰ��R��'98���}��T�6��)�z8��G���%a,�x�~��=��cB(T