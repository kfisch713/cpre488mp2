XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����d��Qw;Z.T��^��P0@���{��`���bt�a�{��#u����f�Xh�{�*/3
�������؉�u�Y_{�@`�u�$��^�F�۴И=��BiIw�i�]R�
k^*o�.ӛ�[��@Lؗ��\n�䖚?WE4k=��(XT7���D�n���8A�k��[���U	�5E�UÚ�l��ܱg�z&3<�/�:7�zz� d����1���'c�h ��V5���Gk��S	�"�H�l%jW~���=��Ү_*��Ԁ�2Y<qM�rX�����\�4#/��<�+f�� �N�?��;װ��CVq5D�H�63��Q[�|Dfct�(	���<(+r����RC"�H�E�wi~�A����m�E;A?��
~y4~8Z�b��� L�xE���A�g���Z�)�� �?�!14څ�?��3�g���1��g�+���{{p�B[�e/C(��,���\?�^.��G>���0���S�6�4zOCx�)��n*�� *-�W�=��Jo*J[w�D�K��`&հ'�٩�x{WpM_[8#A>.�j��:�Z��p�cx5���1�5Z#4��x���{�"ԧ�th�t�d� ���Ɉ����d#ៈ[������c�UOp{iWy�h�̅U.��ld+��#F�]d-���^�"Z=J��.ѧ����k����X�h2��Q
m|�Zh��W0ި/��p�Z�	��81_���ҹ����ա�:3�f�/f÷�p�U��d��
��3��I�XlxVHYEB    15b2     890��ߎ�kd�?�afxeZcC�H�@v��9	(-:�����a0F}wd�*�lh�@!��M�M�ꠓٞ���H�un�B�x������p�(�h�t����s�����G�X黛��6��47iW�GC���0��	Lr��m����`��5o
P&�|x��3]���Xmg��e�s���t��;T|.�j���!Z�bb�/�.OcS3���s��Z������|�b��а�2�H.�r�0Q�J�m<�.��SAa���o�F����F�h���A�eQ�$ʌy<��&�r������������hN��y�˗�x>/J6@"ﾇ�NI�r��5Q�
��˥F�^Y���0��u@�G��:������a�J���k���.i��3�T���o��3��hP�C���?��xJ���`(�猟�hr����
5|�j�n
�{��&�:�\U t<�?;�15�p��N�YK �P�8f1�Ϗ�&6��K�-.���(�)^ˡ�/8eέ7A�VG⽱Of��ywߜ;��a�ه^��]�J�'�˃	��q�X�6wSSX�n������JeLّ5��ςp`͛@`Ԓ�l����*��Ӆ�`I\ �����/P�&�l�T7M	��I���P��l�TkA�_e����Yz��5���~Ne1���V�>38�F�8$�+l:����x����e�����q�����st�QrN�j�����wa��%	��aY�nk�G���}k��P�$�k�G� @r�O�L�y�.���|���L��-�w��g�)��L�y�D�9C��QԠ�lN��jՆ)i=іA���~�g.k��)�g4��ԙXJ���)}�.�s��r�9Wtwi�Ӄ����umc�^��u�*}ݏ9��+�O��]�y;{��l����i�(�`��!џ�'�f��9��R��u�:��'�aa���K�ܼܿ��h7�۷
(@�D.�!����0	zX�l�)�ʔ�����&�)����肈]D5�Q���7�%{�`I�Y���j�h�#�=DW��Yrq�6v���7ѡC����eT�9���?�N�|]�k�oo{B���<����鷲��4��'h�{�*�zbr�����Z�1s�f��?��.E��&� >�<�6�A8pI��8H���[���v�Sf�p��a-3�Pv�7�ף�*$�+���^�f;�c2�Y>XA��Z&��ws~�G���$��vTL�k(�8�rȦ�<т�50�wl��G>�E��������g�(�]���\XV��@>��v5<]ил�e�
?��q����&�J��)�$zF����d����s+��X�_@�k#*mn���n|w�Mfp�7C��{�`:VDX/I�Y1_�D�i#²?;�91���a�8��3I<���觾���_!,^&l#�E;�Hm��h3��6�/�5�[e�J�n�B|�e����9`�nf%{~>�Տ�Ĩ�KA�ɸ=�XVkI���MQHZK�g�+�T#$����WY_j��9��
�d~M�ۗ�$j��	S�P��0�S�=��y�S���.Ks_u�k�y��?�j�3k �������2������h�e��?�7�e%��X0�
������nPJZ(��<���E͠�]� �����oz��/�L-Pux�q�Wk��j��$R������qS��W��K�ح)�p��k�1n�B�G���̽$JP�Oٖ��n�0������~�g���(���q6B�m1k�g�\�Jƺ�bO�s//_b�奍�s��J��C��v�������[�~�8��K��*:sy���эE��}�����x+��i���|,�ADs�D�SCB�$�7�bǷb��\Jw.V6H�D�Y}� �� 9͸InO%��뼼b�h9OaY����N4�iS��%Ό�6g���[�$e�i�?�p��|]�tpdwܭ?W�!�븬6��\�пx*�\9�,�ۓ�<z��FZ�&�W������d3#��.&���?��m�S
��S�����3��ɖ� mF�2&GrTD�67����'^y�����u=k��NW1�Mc����oQ��Y�;��wVH���-�(��@^<��P,�$&��q�����h�Ԩ��9��k�z6p�