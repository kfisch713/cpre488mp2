XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����*>s�|Ϗ�;lE������)��IE�q��}z�9ͽ�+ke���Ɂ5߲q��5�e�������\���^u7ѻ�Dw���:X �|�:�yP�F�'��LnސNDezzζ�5)���J�����8�5
>�='�+�t�������ܵF<����\p��2;�SK�b�~%�m���:��G�!N��~$�"�C�����P=M���8�@T@)�̤��>��z4�>h��G1��Ɔ{(��L�� mG.�"o�FF^�6� �������YKH{`U+Ce��5�F��,�SV&���^�^,��2��B\��(@b�*��LL��vK]��t�m��W��VF��aK�Ȣ�+f���]� �Z��kL*UL{P.���`#2S�b����c]�<x��뤝Y��sٔ	��x�3 V.��*[/���1���-����˼��2i��v��H�ψh��Y��A����)ʇ~d(i���.R��1���Y~����L�P�k�^KўϊV�����7�ƃ����΃���u۩�=0O�]���P�FӸ'B`xz�����{B�;�g
gD`�\u��1��xI���]���X�����'2FG5v��K̄�W����C Z�|�V�nI���,mx(�(6د�s�]��<OЉ�ĝD��"X�q��B3�̰�w�� ݚ�y!9��)�zD���OY�&˕F��p��V�r8�ƤL��aû�)�ѡzk�ƥ�yX#kn.��@ZXlxVHYEB    3e93    10b0�'V6c/��'��Z��Q�����l��V�������e��X0E�y��~��ȡ�o�e�K<�5i<[�܇��A���"����IݍБ�ӎ�`�)�Vҝ��'�E,��6�Dn�mt�%�-�0�g��άK�T���@1������ի"�+�O�I�5ؑ�p�p�iS�t�ϩ�zAyo��# �*>C��&t�s&6��Mxm�~Vw��$�X����f�j������ֺS�<���1G|%g���)�~��ЪN@��b���1������N	��;$\�P�U<���;59�[���lG%�r��2U�"J_�3Wp�ٻ�v;�5Y�U��,q�1m�Ӆ��g9��/�f�YO�}�
|8��m>F@m9�4i*1}5
�h��h���B('Fҥ$��P�W���������F�-�H�4p)Aq`T��5u�`�_��I8]��s�Ss�XH���_�>�,5�����)�nU̐U������jN��V)����ƍ��q�2jt9S��/L��;Q2�XV���8­�"��U��V���N�/�X��[�v� C�:b�hG��;�;)�W��IkpG�X��2��Բ�٤�~�|4�V4c#d�rS;w��+^��3�0:;&�j[A��ֻg��y܈	Q	։��2�o�?3�~�b�q�P-{�D���G�v_x�jmjq*�|Z�F\�'Ѧ2H��F/b�y�zI�wH.�.��`5P���K����M��Қ�}��m�o´�\�.4Y�����sϜR&3x�y@�IF$�s0�=B#�W����߭�������Pn��<����qw�Y�F~���6z��B�I-����r����V&�}1lMߪѧg���h!�4ˌ��P\˔��$7:�g|H9�	Z�=��|g�FO�n�>8G��P�5�g�GWu�z���37�`�͠E3ϛ���Ć�Z˄��	
��d�6zR�ȋ��av��\L��n����y�Ƅ��FmQ���������p���Y�`T;68�5��n���6Jc�A=kWT����{��(�E?�I��5��XP��1G�5f�<���^��:�h꾏@�9�	Zl �X�A�+^�Am��+�]��YR���mC!,"�`��Z��qas�C��hB��/v��C2[`�4j��-���`
�G�Қ8�PIm�˅���x}a�+��"�#��Ih�{�x��ײ���z��N��ø��ɭ�vū�Ȇ/��u��s��46����P��^A���!���x��u�7+澁,:zP{�&Ï������8�:�O��c���
S�X��u�ݳ�Az��T@����)'~?�t���L��r~�FB�8_h�b ى0���x���!���_${<A8�9�[��@���O��d�ZcݍV�b!��M�p`{յ��60ұ�1az��Iɓ��Bf<Fs�P�r�����I�*|e�v���Or���PE�3�rY���#C;'N
�����Q_�o��em
]w�qVz��9�����K�,������X���c������4��iI-�VJ��<�ٕ�|ȗ���>öN�ǎ]vk.X,M{f���h��Q���l�ڱ0�;���n�u�i�J�*�g��[��u��e�MTe㦼��H7jw���u���I����!߫.��I�EM����tJ�GU
�B�����B����|�g�l/�.��u_�Byl����2�>��-a��o�8��t`o�M��f��Q��ϔ�g�g���{�b�E�h�a���>!�Kno1����4�&�/k�*G�U��N��R�c�y3���7�mu�f��T'�e?��Y�b�L��Z��+]Z?ϬFI�F���{��*�ݖsi�.�oy5[��Ml�_z*
6����.wO��/n~z�pC%���O?��k�U��9mf4��8���*��t�F<5�@�0�����/����c�X3[Gt�	6��A>UU��2�1�m!���3;4.��@J]lLz��g?��9M�;d��.�~=cT�9�u�����x6�`m�b���^�#1k�*]���q�2PDF�}��9��"�@&��'���>���~
�rY�oY��U]����=-�	���G��V8Ժ�����`^���U�
N=�����>��D�8�d���±��ƽ z�GB�_1)�ʱ�QYQ��؁|�������3��?%���fc^,,�;݂�9R�n�J�#Xq�ߎ��<�>��1S��(�r�j��$���N��(�WZ��ػ���=�#0S�~b�W̡���垈�6�q���4[�R��_~�LR��+�٬ڕJ��o������ļ��������<k�щ�qQ���j�/jl�����H̒C�o�2�}%b�N�@S�0l��X�	!���+3�A�4��1��=�P I�a�����'Z���2���fxr�K�Cy��i�b�^V����v)-oy��>ib�?�'�;����:bNk��.�W����������d3&��,�CI�<�T,��~�w��*WҬIg��ݏc��38|�]U
,)��}t���6�U�U��Yg��I��4[�/l�*�F�+?����=N��f(;�����;���� 멏�N	�mS����W��7��E�������#.y�"��u�M����m�<��T!����H�����(�Y�̐�c(�ȻA��	�v��]���/q��i��?��y�P8�P�i�p��#H`��ħNa��鉊�"f��YRݳ�#���p��
 ��#�W�So3ѬԎ6��¼/�����Q��E����4A�/�ڪ�;�_&����׏b�Fרa,f�_%��� ���ն�������lA�>��_�.�̈́Y0��N��-9ˆ��`S�����Z���9�p�-��(tP���W��9���|��\s�hBD�?�15;0�)��G�尦�)j�:�����$�Lc��Û;�C?�J6��N��EP-���V�/�@��&~���Qi��Q���7��E�x�����y�1��P>�zg��]K"&�L�:��P�lW�z�I�K����wѫg*�-�O�ں7@ڋ�:zծ:��c�r����F�r����Z9�|8�ҹ�j��;������hD��W)l�au��O��j��j��Q+m^��܅�P�"d]�P����3)c���XJU���wɴ�2��}e���4���B��/,- ���r�{�|&*;	��i��9�d��a��ߐ�
*i��n����Y~<���n����\1:�Pݮ�nG�B�Cx���O��j��>0��GrGO��?:��¬�݋�Ǧ��1�j�Rҕ�(���Ξ���>�s�A�U�P�bL��:���A�ID�?�}�Џ�_�ʳ���!_m���a��&lEM��Gc�M��pf�9O��� "��pUC�U��w�c��'c�׈�z�"Lx��⸿r��ej�&��fnǁ����~��Ê�s��h9v\}\4�-�@5�����@WWɢs@mK��X���ĥ�?B����
.P��&�=���D�>,��G�
f�J��G�����<긴Ye���� �� PUK!�(���M��� tK��:O[�#��p(��N�k�L!ˎ����Ry��y㫿e��}���Z������of0^-@���]��F+�&�C7��F[�������*/1�>r-���9���	f�a�t�w�ؓ��3F(�mڋP)����{��ۧ��UL�7����y��8��/>N�ͪ��� �9s_�O&蹇�� ��Q��]�)t����u�����1�-�7��a��}��i�0��o�y���k��v�'K���z�%�J|vv���Vb��F3�Ri�j��ˆ��Tڥ���Q��"�D�{w�J��W)����eP�����|�Ҫ��IL`�}�"?�hkV��K	#���s�+�V�ƛSU��(�&�����	H�ѕ����4WSeq�x�48�J����ͺ�`U�������It��F���<��d4S"'�So�~%D6�a�G3� ���4{z����}p94D$��B�H���r��$��00�g\�hWN�u��w��d�.��L�j���m����qNh�r4ȼ:���Ec�b0�]Pl��{t������v�(31�����)%=,͑���	����&�62x1�ܺ��p{>��