XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��⽟GPYIY��*��/���%�&*X���7H�9�Z�2#2��9��gL�� 6(-�ʉw|9�̽�z�B�}�1�<��׫������JQ��Z�A��n�8�!�C�z�RJƴ)�B^���}X����ϐ����cpR8e5�DU-�� �f�A�.��W(ʜ��A�� dc��`.X� ��:�`�$D��6��޷� pE����c�I��gQK�RV���L�Ԯ��	,[��3|��>��ݥ)Qؕ�[����~����#0���Ia��u�7	<��;T���ߧ�5�}��".�-�o99���[?[i�JKg���Wa�'mn����L������G��t�䯼~	�dS�k�O[be�b�jL�$���aM���as��/���� �
��|k��&��r�;����`�5< �X{!!2d=9�'�3Ė����:'�{L���3T�;q8��Ga`lG��u�o�d[��Ө�Y�|��-*=S�`w��O�͒�V��
��p���[��xa��]��F�ALE�y�P�(�ݶ�u�F��DS����Y�%�Q��,U͙�$�_�V'�&���pA�dg��A�n����,`��o5�c����m�	5Ԗ�mݠ?��8������Ƥ+��il�������C�q$�R�}P��~���!P�|
�#��"������$��uT,;{���쌩A����m<�};�,0T�w���<0Q\���Dy一{q)t�fq)j����_�R��LXlxVHYEB    b087    2540��a��{�)��^E��.�Ӌ�_�poWy�o��*Q�>: 7������0?�s�-�v�=�>x�I�~�ILJ,h�u,4�i�W?2�d�5Tj��/.���:�����.�W���痦V0[?l�c���R3�Dݲ��Ju80����N���^+�hd�q"AI���~�R�h�Qvr�d1�M@����x�X��-U"شmdש��L�O��|z�\� �a��{K��h7���w�����(�ַ(�0��@R8��1a�'l�G|40��dAo@-�
�3��C�Y�l��Qװ�EOz;�m?�����L��?����+�ha��f".� :/u5���Q;H��P�07�� ɵbc�0�aH ��4s�=s�]k��~
���3W/@I)M������IF'���q	�������r���rh�Z�J�YJ�D��Z�7�f��Ne�ij�-g.��큹7�ߗ�)RG#�r~I�ؾH@����j/"T�#�j�Sۙ�Hr�J��s7q����3����րA�G�'�ۇ1'{�p.X�Jv]��Q�6�,g�E0�4g�{>x{��M���R���M�I��C�� ��>d�(4+�SH�����h��Dj����P�Z%���\:"ʙ�R��D����,�J?��S����N���3^�X�ZjƇ��c�q����F��j�ZԮ���οf����C�����ܙM�p*U��.�0�_4Yyq���"�9j���W�p%]G�f�1��p�'�F�u���k]�������m�ʧ҄��t!�Ÿ�+Mq�(�=W�ìq�@ȕ#940� փ/D���\��L���)�uw]��ow�1�޾������m�n0��W�����f8�ʰ��(ծ����5q����OF#�S�l �!��Ǒݦ]o��UH��`�� ��pEVfͪS�(9!�����V?4�>�|�c�"�8(�[�xe�nc~����P�e�o�s	�n��i7�ȝ�y�dJ��
��̃8��{z ��ژ�!M5#P�6xz�%Q�>��3D�#(R#8 �ߥ���K�`����ٽ�A�}HG�"����;߆� �/m�-�# <O�+z� �:�rXl�+��~��S"4&�cmO$LhM�[*�ۙ�K�>q&kl�MZ�����+��a�i'Q|Q��ɷ�Է�\a+�'�4��&HHʐl;d�(�;٤'RI5�A7�K=�<�L�h?�R�X����ɹM��H�M��1븆�������@:L�t� �>sxN�^mY �@�	�&�h����ӗ$�l��Āt��O��Q2�}�`�l��9���� C�,��"`�j �Ä��ĺ���0�]H��*���j��>�w�5i|F3,1{�4[Yɧ��.�����Q�
�ȕ;���/��*QH&6?|�@�O�G�]������r�d���9ט;:{�V�5c�m<���&`a�]�auL#�f0o�
�";�}���­qvm��Gd�2�b}���u�֚;���Y%&�w�o��C%��t�kA�{5�.2�S�>Eȃ�pk�P;+d�x��6�!�)�[b��Ϊډ3�I5Cg�Q4��ı�4wӨˤ|�a�eH^���D�NGGEÏ�e�t�C�(�e�5�s�����6��E�҈�n���J��wE���M����i�G��o�4�J��6��띻)�2��0���j}���qo�>���ʌ����0�+�}}�_��O���-))ف�Aptٚ�.�"�������.Dy�f��"�lǋD���r0ƽk?�ə�}t��5�FTi�Y�~�Z�L���-Bn��{J�����U��J�����d|J%�N:�1��U���n��'��w��l�vt�r�|�L�ЂGv���ݒJ��Uy�?@�H�,�xi���#� @ Y(��#q��CU���^������cY�"�,��p����B�Nl[3��J#��ѷ�����SĊ��Ƹ�h�$!�_���a`�c#q9�9���j��5p!���[HI*H�=��#���K/2s{�<r�y
a�r(�3=)�
6fpÙ� ���������܏�� ��"�rm�MX���j��3t�����en:�,W���(�=]�ո�h�՛`����h�O$��3��o�[��炿~wh�|���<�K�D�f��hC>i�q���lc��c�-��S���������g���h	����|��y?��D׋M��?����fv�xo�%���ࡿ=v��k?�,��E]bF�(��#[�T��⋿q#P��*���ϻ��sO�=��P=�_��"� Q&�"�Μ���_��&ch���]���O*z��2ך2Cp:z���	����R��a�F̓'T��<�l]�[�UBEU�py�6;�k�C[m���ZO ��,�Jl*Z������jO��bg�%�<�Z��P3����SI1�[�z�&ϒeF�TUD�P��K�cZ�0��]�8+Z0 �>וno��Qq �)�D��&߹�1x����wBE=z7?��Zac�,*X��g۸�pjp_�)��2�ZtH�4�5��Fv�ǪQ��j۲}�32S�H��m@+UJ91>�'*�먴d.�'[���B�oo�mz�����-yʙ��aN�Z����={�a�K	J�2�o�. ���ɂ�lW�i�֒�Z�ZO,=�%��6eo������*��/�����}`�Z�ș�����.%�bp����ŝS@)����U�T�I��6��	!od��$��6W�E�i�ӿPq��km4����v6����sYh�>L{�߇� ��[�K&�����'t���jL�!��hY˞�1@�A���,_ =�R�P�ޟJ��:&O������7$�"
���1b0~H�oK!+�,$���x�",_::Mz��_&]{�
t��\�Z��{�r
�y���
��(%�=����%:��
��Z�`�E�u��A��l��]+��]��R��G&k��\8n)��JȺ
��R=n��Ц��\G�Gz���*l�@؍�Aq�\}Ip���Z"Qq�������{2:}qC���,YjF�����-C�f;��͵*�.踉���:�*sG��|�]G��W9�A�4o����0�˥�L���Q^�'$ldRq;�b'��uYo���V�h����݊a9C@����A��?��'�#�?mYP��3�?�Uq�ܑ@��Ǔ��0�o�/����(n�_W��6x��9p)n����=��%Hݝ��}�#��X('���L��)k���zv9rS�N<0h���Ư� ��U�$�y�s���oV����E�9�8Y��5ǻ{E6�Eq�v��Ʊ�����*&V�.�u0Ҷ9�׈�y��c�sY�s�qA�귝I��e7M�4_U6��z�T��f�\�X�G.��"��۠�><�gͥ�[�%���'c�ja=���d�n(Y4���U23*��o1�Jo�avh^n�,K?�&��������-G���o	�w����9����?xl�ʬ�SV�"c�fz,Ɖpُ?�d����T���x���Vz����g��27y`���a����_���{�[ɤP�]&�\��i��>W:rp?��I�=��B�FU4JI�&3��8ʁ9ƀ���m/�F��n�Wޣn���__1 ��+�l���J�<�l�C����|�-��?��u�P�n-`����Zd��e3��`_<�$�B������2|�'p��I\S�
�K�d��A�Dt�����zO�҂����=��.�M��o*�&�h����l�����$aS^}��/&>���T�M#�� lTc��M]L�����J�]��t%ġ����߆��4�Æ����j�4'��� �Li�ʼ�>.�����
>�wY��J���&x뉾��*����1�#���U�k��ؖw�/��b�Ѥ]a��ڇ-y�B`��;CpR!��{��h���-��B �Ĝ�W,��m%��HIlupO1^�J�����9\�%I~���7/C?��l�ZF���`
"T`���-����&T �X�$��<�׸�n'��lLH�Y5�U>X]x_D5J�&	�u��)��7����f.�
.V�#'C��ڷ�J��Sl%m��*�Gf����h^��F����qdz�2⟨$�[��b ^���#,j`�n�{[|Y�Y�� |�.�������X���<_!�`(��xQZ�_gT��x�:"�Ӏ�1;čq����5��gV�T���$�����$��u��ej�7�Š>��y��f�l
,�c���"��>�n��1��.������D���gzfMW�e���@^q���Aљ+"�s�(5�y~�Щ�S0g�$̕����c���w/�-1���/n���p��s���L��:��>��8�;�5Y�8]�Xia�(�fA�&��Z�2DU�0�h��+��ɫ+���HJ��*e����?�8��zZ%1N�B#nim��]�QS��s�r����� �?Y�b�`�"h��X���\j�q&%Jv��!��k�|=a�/܆@Y�a��ާ�&�� '��p�W��J����G��ث��J��ra��3��5	'ߌE�;D���$0�X��Tx@6��O�Ö�S+2xG��*��!�Ug�P���Cc�,@(z���<<�
SV����lY|ǋ�+!��Qi�f��2&̘�I,1�K��������=݀ϴ�`�qH��jI��,�c$�㻢�
�"t63���t���*>`��9�.�,ؖo��|�/�y�Jk�m��Pm'J'^���|s�y�Y�=I�����B�ڞ?w,[Q�(ք��U^��H�A�1u����9�� #᩺&E��rRt�Փ��Iy������̕V��$K�' �z�M=Ų'רi~]��~��7��Yǯ��$A���}Ea��o��} �L޿�$��?�D{.ͥ�ч�B
M[AtI�ң���;�����pEV�긌���h��=�'fr���?W�e�ޓ���Ջ��Dy�ct�~�gf�^ʜ Z4IĒ�Y�7���ps�U��^��:Nϧؽ�]E�o�dm�yVk�~]ST�!�/��^U!�+��Q�V���i2��9�u�%���Yx�`�|;dnI�_�hmB����⪫;�4oM;qO�jd#y�s�_���"T� 0�����<:Q0����V���>��(y�P��ϲح���m�>�O���Au��g`��8�?^[��-�4�{������(��djJ�0 B�ĨA��Wq�vS6�,!�%!Ɖ8���\<x���YI�ӦMI��Wh�~��]ە9wNȩAq
�7	���#�#1�*4���!R�^6�Y���wRS��������G����gU 튔�	���4T|����FNd��#JaP��~�f�.����Ӑ�5�?� ��+eBmZ�)]�����,�g�L�3A�1�0F���l�s��o��t�la-=^���1	�x�s�Q�W*�#���%�˩��g�T�������{m�+���rC�j2�� K�7jU4����D�% _��2�7Qj*�Q�V���4��� ��`:>�h���nU���%��Wn�>1�)̭%��D	q��n���^*��љLa�r1J\�����3f��J�`��I@���J_��x�8aj�_�����oS�ŧ����so/UUr!y���]��.O���$lM8B����)��t��۩ʎh@��6�e��Ku���o�}�;�(�`[j^[R��f&�m����'@Ni��]L'���&��	.,o�R\ ��!AZ�^���`3�y�ј{�ŧ�As�����F���zz�Pޡ���H� ݿ;�[V'�8�J_٘�mr!��h]���Yq����5-���؝s;�ʒZ�Z���� �&w0M�z���[?�.�I�:���6��x� jn+�G���L�??��\�_����y'ψ�"2vጓY�?w�kz1�v�G�D�a�g�����(U�g���:Vs�f�ʽuF��Ki���躺��L�3���r�s	6��t��Z����.��h0���ٶhR�Ί�	��#��L�H6�pT�W�UϬ�)�y��yfX����ශ�|�C,׏�"Ɉ���M§+��8d
���6��V��#��I����0�j����v�78\���V���	�ĭd��j�_ę�x�H�+�
L��p��DL��8!�����iTe��t)���$�J&Zط�!� Ts�|.����{��LZ��&�|�1�zے9�=�ڈg���}�+�xi=��N��h}�2>x@�M���k��]Wv��k���T�y����
mr����_%M#p�������&�����n�C��@q%����]+�{v�(������n-�^@��%�`6�KŠ#�1����k���p�qn�}��׬Iբ��y��&����D|�R���92W��{���}����������~����=UP��PGhQ~=�8�)�2hs݁�[dƁ�jiTAU�ަ��z	�o�N��`�.�r�2��&��($}egb8:X� ��4$k�A��`#-K�U+7��*�z/&��Y�����q�|�й�k��JPE-v�!��wqY�M�!��}�oX��<8�q�Df��j��G��Gr��Uf�@"٬��n�f�*o�ƇB!:\�:e��n��Ԟ|��!BM76���{�!���-Z�`��sI5��3��])ٌ��+^�*b���h{SXH�E�o6���<�/Qj��;�6\�>C}jV/r�0����؊6�Ҏ� r�`�T��Vh�����p5ˮk�ĩ+PMM<�b�1	�s<}���ân0# oL�N3�V�!k}mM�DK��Yj�p�8/�T�M�}+�(��)sK�	F�i���9&/ɹ� 2�2t�? ��&��3�pz�.�}y6etѩk�DЙat+9Z pl$�p�D�V�K�ة���o�*��g#�&��e2�bzR,[�*��_ۗ�4�/(�x�42||;G��ԃ�QF9��wg�O-bG�X��T��bT�G�`�zD���o5}lT�eϧ���*�i�-C'�"��c��F[�X���?��̍V��Wy����՗����E�-m�VY�BR^U�~��Y���4-�6�6�Pj5��vܰS���p]��^�!$��vm����Ohl�^�]ʖv/<8F�n��H���2�gn�.��A�J�^�(4	��\� ZQ��OK��W>�y]��Ι��vad��P� r'�)�Ŀ���0�/sڽ�T����0b$�?�������*\%nw3Hϱj�_X�F�0NZ�z��]W1Zx�P�I����{K�Z7'ч��c��P"}z�
�%��]`��_O* H|o�A�B����.��7�ML榽[4W�)~���7��Z�*��2`lZ�[KdB���?��?8܏j�M��� XZPR��ȡDX�~r,�>���q��%��<��yN^��q���hp(�(�!�DS�sn��a�>���x7^*AH���Җ�w�6Ii���x�b��uȆ��ᇬ�W��`���h���G �ȋ[����"pz�d�1I���8��$p"�1����}8��}�N=���{���S��-秂�j=�mf",eQB�ֹ,6�IP�7�Fr�a����ݰ�ƴ���X���?{� ��a���U�bÄ64z<`&j"d5��-�64!KD�Y���84�d ?o��Nd^��OI|6:�3'�����r$w�4��,��q�`��Ͽ������T@F�����_����,z]*4�HJK9�ӏ��آ�'{}�����y���c^B������!pNx@��m1��YR_�h�L��>�.4ьi4�.�ꄅ^_>f�	����nV��s����`cʛ��v`���xG�8���I�}�"@��"�nAҼ�ql]�2� ���r�e�ĐH%��!�g�m~+xc*�P�k�����MP����}d�����+�/�z���=������wn�s.��CM����?2�-u@���K0^�b��7U���D|}vU���R�5K�A-a�]�dM�%�'"Z(9�
.0���ߌ�p'\4֬N�V^���х)^�l�G���k{4��$c�2#j=�aQ�$�b�?R9��w�����b�re��G(9�.���VqY��Wnf�j�q��P�J�Z<b��g>�6�<=&F����؄#�?[�ǖqC<Y{f�8@41�(4 ��k�ĠS�0q�З���jYO��wI87��'d��f�5`A��%���IM\K�E�G)���0�c�����7�� '�Rm��mGę s�Dv�
�>�K!kX�靃�n��K�@��}6��GN�¹�e)��\��>����(���S�}a��	Dd�H(�7
Dh������{5?��t���2F�f�j�������F�{R|��կo�#%�\�:�x(���N#X�����M/����� �yV�[�u��"M&%d�f}��cT7��0�~��w��_ek��{6�Z�"����o6��i2(���T�IG�����G J�l�̏:�q����>\����΀�o�CnIv�ko2��y��}����Z��%"�K����Gt�l�MѯSC�A��mwa��\�y���pA�)�枋�q��= @�
h�	�uQ��0;n�_��.�F�#�ڏ�N0��:�x.��oD���Af�z�p�[�`Lwu�� ` 3���x��M��2���θ�u�#L3���QbR�{e,ҵ��XT�/{'�o�]%�����qd��1�՟m�����.����~"�`�[��d�f�n��_��������W�!mC�F���r1
�0����8ݧ�<#�]$L��I�,����8ص\��l�v
jۀ� ��݋\\���	Yӂx~}�Nm�
e"eS'�1���a�>�����}��pe�BO���3.l�%Ў���l�P��b��?j�X��\�7ۣ���H.�Ë�<��&���p+!�v� �hYK�4���*����C���&d�;~�'�-�A���{�����J����_������-��ro�P���;�}�t�A���N���&L�v+,��Y�S����6�V;uKx�ǑM�c�"�)ϛzX�>�K�3@��z�F�z��O�sG��y7k�7��۩��!s����]"f9w�za&�.]}BO��T}k}EH�B(��c,J�����u��;헅�V,�hlv�W�g��聆X����5\'����D45m(��ā���x�J���^ i�ߵ��Z�s�
(I�|?%��թp-�
��e�0��L�"9n��4��u����1����b/ļ���F���y1�E�So���#��~!amr[��8ng��YC;�gp��1��-9��C�{3w�