XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w��߰v�C�1{D�8�� ��{"��D~ғY�F�֒�r����&���U���d' ����W:ޞ_/k��Mkq?�o72\ç������}IC��K�F
fj'1�P��/9r�������.�1�,����u���_6��M�>F&�c��VQ����������h��[��������r��Nm�8��~���Eu�	ϸ�4�ث� [�Y�Eoi�I�S�@���2-F�B^�%F �1\�A���,H�W~���fc��Ds���,^��?�V�0q0��̘�� {ީ�9�.��&�6��!)M6�ܳ�KJ����⺎.�tk�:�G-�Q��DYclqk\��i:�
nWT�4���Õf�iQ�S�aNQVy�<�ގ6�%� ����>:�V�VU�+�p�l���ކH��!�����Q�(xfs[Y��	��v����x�>5��Y�o*<I��3��HS�۔+/�@�L	I0�������j�e��	��M�]�G�eyg�t�Qh�
�a�Ze��_�H��\Qa9��m�*|�%tжB��������3&��T	:�n4m.%�ȍe;A4Q0;�'����0[D~Gj�`f��׸e����."��˂Bz���ƺ�\�#���:�Gk�e3�Xv	ˁ���`v6kÆl�s�sZ=�s��[x��x�G�n��4�c�Ӄ�\��H��	��~V^�7��{�#����͌U��C�a�ʅ��f�(���h��S�c&��lq������]��XlxVHYEB    9fc7    1fd0�����#��*/�l�"��^ۛ�����D{�$��y� �\e&v�<,��'�h�[:Ne�Hx�ٺa�{b :�8h��ʋ1�2B��M�i,O�=Ŕd.���h$��׊��ϛ0S��P� {G��P��W�� g�P,+�>�'s��-���Lo�T6d�"��Io�y��`Ez�n|cv]���eI��HqE
Z�g�GGIH�m/*�G�MB��r/���2HX��E�DC�B�ܸ���?��d�Y!|����Ǆ�\�"xh��AX���`<��hԚ;Ir§�X�2 S�9jB<�����,�I�(ּ~w�c�x���;�"�<���*���9L�yÌ`�^y �5?{taF�B�tS�'�d.K�Z�k^D�W|V��7��Wi<��.:�)R�,6����Z! q�,丹�~h�?cSZ�Is%��̜��E�`���8�/T�k�%��q͘$���0�U�%������Sǫ�g/���(�O9E<�..�c���'�*��8k����A�ZI�N���@���:tp�m���]�? >dv�Id{=�y0l���-6���E�
�b쒣r ��	Q��,��A(��^��C��E��i�c����۰��>vwAw`/2�Msi�ίX�T,W�u =�ФBx��BK�Ǆ����UM_��6�BT�i�ݬ�$��!��ФF�y#Bxϖn7�v~gśeh ޭ�u(����%x(��l:&�<�q�I��{hu|�9����]^.�/My�vk�O;����@4l�;D{A��ěk3l�-]�eTh��b��F�	�K�cn;�zFs��}��>����d���uO�YG*��"���h� q$��H� ���\O,��=�<���׽��7�{|B�/t{w�#v�7��O%�Xg�|�VU��PI���:p�&���^���%�Xg>�|��A���F罱j�(ee`���Ŀ�i��ɢ�sF�V v���J�����8r� �����YK��{�b��R�Fy�*w�}��'`��S���v~��>tP{��&�|�jd�nɹa�64���^TOx��0"ac�ST8�>�hy��}W��C��l&��ʪ��ϔ�x3�T�7�5��s��U���%�xաS@T��JD
	"��:�l�}�>�/��O��<�(Ձu=!��<zR��>P��ޥL�2�/��x{|�[CxI��?�T*؆h.I����s7]{^:@�� 9�cGq�8�$���}Cc�h��{ΰFN7�	������S'u�q���pc6��'�5p�ek+b~�2��L�P�h����j��؎Eo$w�˘��c�6~���ֿ�ĔiA�i}Tl$tu[��K%�ػ�X��?:��3�do��څ�+zX�����R�b
ç�ܬ�c���MJ���{�l�º�q"�AEE�i����X�n��t�]���r���yD���)x`�@sښ1�1;wⳄ�g����(�7�[(���i_���S���w� �>�Z��̏ ��t�!Q���@�ЋlA4�G��sq���Re��^i��$o��=G)D�C:�p}��7�+1`}'o��l}_4;�k̙� �WS���j;�jIqL��z��A���:^��1צ{�{L�D5'f��P��ZgQ���oM����MI+Aզ���S�QK���w
Y��;>��XSA�y�M�{$�h�]� ��߂�Ł�)Dv�p�[/�����C<-<�H�dB��fEE��a��,�d��\���%2+��U�2��R)�K�"�*N�b�(�9�x�i��k卙��;�r	{�f�Ӎϱk*�-�N&�Ů�w
	/ Os�8a�}�;�z�P��=��$���)uv�7/�S��M�$��(�g�g���@��<��uC�P�I��pnL;10S���<�=V{���:_�|�ΤP�L�.�}�tC6_��z0̮��>�P-WR̥>��6�?O��<v
���R"G�[����}U�i30��~�3�q�W/]��P}���;v�k=?�X���T=8�R�$gIVoq�xb��$�}p�����Ze���pg�-����i(oy]i��F�e����H���)]]�N
z��T�Wu��[3u1���+��X�F8�7�xձ�~(�խ�����G�V�n�*ďy��
���7d�$�dl9C�wk �����S�K�$65�a��(�ˌ��c����,�+�;/�U��_�y�>�����9.��=���{�\ql& �"Bp�(h�y�I-����2��q���\a������Z!u�}-�2��Wl���p8���%�
8�g�쳾�fa���U�8M��H�����^�aׅ �'-G����ඐ�Q���1 '}r���H'�8b�I91�u��O�OP9gW�<�=�����m����aԋ��ԭ��w�cLe7��0�]��'1#e���\<���/�q�U\"���度�Ϯ~����Ff���I5o�� s}#����>�+�(�J9O��I��Ø.�j��g��lh��+r~F�����f ��	's��M�������~�މAƀ�v{����5�>۾�}70�qO|	�,9��/�J�>m� ��AR��)	���K[P��iT]�_O#(Q�o8,$ߢ�×�;����G#�6)�<C��P$����jWJZީܕ+*!g�r���K�KbX��)"YMÕ�[~x�ZW���UBe!������,�`C���0������H)�).��+Z���-�õ%D�c��!�F��C��b�9�$hB0���E�����c<��aZ�m9u:��8�g�;����$�)/G���΀��o�09�u.����畼G鎃���<�q�oQ���ykn���J��.�?l����6�̗��>�GL�+0,*�T��\�>���s��sY�l��9��)a�j����qy/��4m&��n�[U��6�Lis�D4���%�'v� �T��YN< �1 �2���
�q{�:�LQg��/�E�Z��2^�	Ve�};�8�Xem
R^��k0wGȅe�E��	�iLe-"=Q|a���(.\iy�)���rIԉ��nY��eq�g;/FV��}��Đ��_�����Ev�Cx�ăYkyY��2F��9xN������Yj|���%.fg�}�.0c�Q>o�	��`�mj�~��>� j��{���\G�y��թm˻�RcNOxZ�Q�V^�M{��V�q|��=xp�S@��ӠrwB�1e��c�s]��W��: �MJy��ż�^h�y4�Ū=ֲ�a����y�.]%�k�@0 &�2�ܾ����:���*lnd�b �:O����xh,��?��65��G�d��J� �������� �XD����	�(��M�*�_��ba:��I�cR�MVF������J�>��Fy��|��K۶�z�x�Li�ݚ��|�_$q��&�Z���ra���YRBx���qm�
�l�4_��ɳ�^�H�����tW��*�U��v�����3%+�&�?W���_�g"2rN�1��Zڮ�rܷ`��z&� l�z��8�����Q�i�J@f��n����hcү��6�"�����F�N�A�w�zgG0�b�F��Q�@��6�qv�l��6�Z{ٿ����Զ7���#h���Lp�Zcg�8v�,O�0'Y9���2�vP}����R�b�H!v-_�f��$F+�z1�`OVI�k �u}�]��fX -���j����ޱ�J.+��$�&d���g�79Uԑ�^�|����w�\�k��Y��#�m	s�)K�.b0f����C՛�Ɗ�R�s�Ao�{��e�I���?[]��ͱ&�eo�bT��b�#�=��((jvە��Y"�&ۯ[�M�1
p����~ ǓŀS�/gw��� �4����|+�@��8�% �S��5@�梐!��P���Z�q���.=���[�AH1v��^�����y��V��Ù�~[�z�bG��J e�.!�Ք�j:�)�[t���~���Un�sg�Q�X�V#6�$h��\L��[�/+�`ƀ?U�u�ZF� i^��^sb��5Z�D�Ѱo�ҽ6���M+%#K?8�a�r�QF�>�ߤ*VWxϟ���,�[�*;��ZaO�����!��fqO��
&7\%��4��f�x���ht]�����Q=����oP�yE
s�ic�MZ7�y�Π4�(�����
��3S�?G��5��2�=�D��5p:�T�`8�%��������/����~|�KB߮�sތ�Z<��)���	�d�R*�P�Y-/���R$dd�n��,�j�8fQ��=qġ�؄�X�0G�reU�'.��84/��:�ҼP��d�mL�]��C���ټ�1~�Շ��쒎�M�����%��	��[��x��<���Q�0��|Q���z�� �͑Ċ7emV���z=�D��I������&O"w 1�pC�-�h�)��ۂH�(���"y�����1dR��wL4$̝��0p�4h�e'�K>d�{��n��N�=Q����
�E�L������z��+b�'�Qsn&!�&�N�Ĝ��U�s�z��L�:���,��/��"�K81u�QZ��S���t`�)��\��Oe���УӄT�HM��E�Bq�i��`�P&�M��=48�������vغ��}�pڰ|D��I�e�c)�(�kds����5�q�G�2�/�;���	���_�zg_ƌyF��)`"��a@��;�5�e! U��D��#��)�J��_b�F�xa_��/�B-��A�0����<>�5Mt��7��IdA�um�8/�΂�$S&-����$B�xX����2�]���޿*T��&{%U����u0�4����!?4꽅��.�������Y���\��b��P�ݚtt+GN�ȉ�0�J��!HL��c��>ύ�d��^�,��'���sA�W�c�(8t����Y���̠�����r�(��"�0i�	 g�tl��X�dc��@o�y��-g�b�:�$�]�
i�o]�h�T�Q}$$cnҭ���m����X�_�����m�tUej�`��s�G*�w8l��[�f|��d!�;��q���ҹ_�SS�B�-e��[�8�Z����������w��V���\��h(pH�V%�XtO��`5��t4����������^���)�j_BȂ�6=�݊m $�L+�ȗ�wO]�I�
��iȷv8y���*�L�Η:P��N������0����:�J*��5�wn��-�B:����!�ל#iUp@&k����QUYMb�ϴ�M�K?1��U6d�_�I��o��g��(p�(���}�T?W=�X0�uG�@=��U�%3���[�4��`�e(���D;a��AY�{GaHǙ�M���tk��^ Ev�5o�ĝ��S��iNb�dyF�C-�x6��8K�g���>���C̾|��,�guR���p�	��A��$��8�}�Lx��4�u�q���k��^i��31��Z���я����/B��q���TO�>	��hj>��Kܫ����n�$���|Apo��Z{m	.|���g/�޺Qti��e�r�KQ��#_�����53�_!ՙ�ֺ�b<+��~<m������k�{w�����>�.N�{,�^�4�aXA���������O�	�9#����K�βVlZ�_����U��{Hਂ�����=״�{�� C�ԅ�2��h5���g����K�06"b��j�c{kc@��8dt b����g/E <%�v���K�"�@FvS�O�T�8��)�ҥ[|m�x�fb�0�:<{�iuzY���V+�7��b+��^��)�NUb�5��!f[�c#9�# ~�,y���ZjA���8;�P>j���j�o^�Z�GW?�kE�&�xQ�áU"�ho�2Z���D6�W y �$W��A!P�׭�w,�Ht��0��S_k�-çZn6���YP�Zc����aS��O {
|�Y!�
�o���z����{������P/q�wW�F[e�qCq3�];v� ���.�H��l��f��vr��ET	��M��V��QZQt�~ �����Ő���ZO�|��uU*�_-�v�ݓ@�x�d�]�PLVgp��$}p���ո�4;��Ԕ�[;I�&5'�þɴC�B~h	 R��[�6�u�ӧ�C�]q�8q��T�t|=�����~y`#Z]�QM`~?rg��,�v3��(��5��ձ~�б�y�a�O��R"*CV@`Lb����,��7_��n 
��g�ZcH�ܰ�ϙ��'��4lQ�:/�`���qvH.��L�6o&��#x`�9|���64��xB��  �1GKp4��M��D��K�/p��#���!��C�+d�~c�U�L8��'��It��]6n��
*$�Xr8uk��>�	ۈD'��G��p��Зf���E3_�<� X%��E��`R�̃��_�4��9Ro��Ó2i"�1{��Iފ�$����1�@[����&�Ҋ�� �x���.�Bp2+���AF���P�u����dLB�j��o��1p5�0�|$�M�U��1�(�����;���M�~E�t��������#s׿���k�Dx�L��`
O�s�����a(�OyXj+$���#�������cmq׶r�y�~E��&�F{��c4²��J��!$���]�<h����4}F�_��n5��{��Һ>ހ�"S����G�ͬ��&)A-U��Oޣ�}��;�]OO���2�.�������R��ǖ*�_��<skD�*A�����9�?B� ���� �(;>;7@���8���|��EY���n!6
)�.��W���0�����n�ܦ�޸�P���WfIOu|�!kQ��Ġ	}���3l���u�'k��H]j�����ѰSj���I6��*�G	���L�7�K?�3ϒ��2���T ��:�#�_���]d�T|S�U�	���N˺9f�jқ� �f�����=��o��Xۨ`_�z7����b`�A7�����׎�(L��g�E<�)�@~����_�Aw�3�i���URÕ"���D纇{X�{_,6'���/�W<�sS�@F"`��5[o�JKs������ݢ��8	I6]��]��e�i:�W���_�K���?����<���=u��(`�sd�U��?�{��9��n�ȜaX%��F6�&��;���5�?��\\�����{O��zc`�Az�@��'��`��99��� �9�RQK�J�C�s�	T�a4����H��
=��)7���tG����)�s.�-߮�}���-�U��7)^�6�q�������!���
h�#J���1�m�r���p)�n�.�=ƭN����IQ?��,d9�����Y�K%^q��Xz���%(ӈߖŦ�������������ΌO��뫑��6H��5l��|��d&Z��I�0�Èu��.!�X��F��a��u��t����\�$��{��e[&��{��L�%4����bG����~E�d��r32��_o&v�`'����	�3JQt3NA׭����:]s�����_�K�ia��h�(�2��@Fg}�¸���:�V"⎤�)�՚0�U��*���F1a�y�$�]c�	�TuN�*�4�-��N���τ�"�ׯ��Ny]��1M�2�FS�r��6���q�@N����o
l�1Bm��>R��A���&D��������J�0�re�z�����,U�U��]=�\�J���`��2,r׏ۭy�"��_O�Z���}4ׁ�f��DH��*?9j����5q��{EP�_�T�g���(u{G� hqP�'g.�����Kv�Q&[�C�C�Z��0���9���h��|�r�j��o�JdB5���J;k���w��`5�v���Ⱦ��Ě���_24�F�`sB�L�+L��"��H��xP�ی�	�d.�C�vA�)�3N�]v:Ch&�r