XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����fw�Aߝl7�H��5��Qcߴ�4�IVt{�`3ʌY�v_�+��b��C�a� k��t�z��FH����'@��}�dq�K��Ҥw&��\�p�^�Tީ2"�^$.b�� �3D>+��Zm`�L��ar�32��3�ue�V�{�F k�[df򥕆z ��_8,,&.%`�L_)��cW�oΚ�5��=��y����78�8cl�)�Ҍ0�g-ɤ����(i�����0��ᬫ�Jk�O�{+�s�nW�[=��{�Q8��dm�n?��.'�y"Ln��e ��:�7���Tu[�^m�Qzb��Fp�c����c���������f��?d�����pLSF1�>�GF-��G���<>'8�Zq�h	��8�oU1+J�m: t'7gcV�>���S�֤N�!o�X�_!���龁#���w����;N�o�_Ir�~���LH�7~{�<O��µLLSs�u����z���k����8��O,o�k�U=)�寠���V�qu~+P#��8�-畱�{�-g�k���w�=E�����F�?ī� Xf��[t)��}�uu���C7u@��'�@K8|/���B���|��=��4x@T�$�~�'x�cf�Y�D��ʤ�Ď
�Q����h�c�!����>��]����>n� x�S�^�0�
��P1ܤ��m��Ǯ��P�-1�*�U�47C���s=��^�#
�z��ޖ�M�M��̗��l��6n�O��9\C )�j��p�Ā�#�V�XlxVHYEB    39de    1170Z����K ��(3�r!$J���yZS�@��|��2IR���Oo���.W�:�%���'	.͜6>Xx���"��2�B��S��>���лް�%����/ �!Ǉ��˚�����(�Q���x�-�������so���3�ٓ%�g�o�2I$������<�T����冋��^����t�%�M��d)�]A�G!��|SS�.˚.���ԛ���E��hID����2��A�a	��~�	����4�z��kW[&�������<;��+���æ�S��Q�B������H��2���N&�����|��7��@���ձҍ����/��.�A�}�~�C�XF0��ͫ�9`nߪ���g���\хl���L>>?�XW�[��$���5��������M�85�K���0D|LR,�؎ ��F�[��4�=�>�?��nu�۫�3�It*DUbW��˥<�K,�s����B����#�r��x,�,Au��F{���2$`�5ɡ�)��F���F��p�{���ۜ��]�3d�0|�(�K27�E@�W�����-y&�k#�*/*�g?��R(?���t~�!�q�(Lh�I��O��o�,8�MF�0vAq#��`-��,��u�-������h��"��"��� �K0��5�*��]���d(u���{˕�}F&"�����yqݲD�G���U#5R*�ߌ2J	���H�J�0%
Zf��ی�W~^"��d������EG�]���?��z�j4��Y�6�s���=E��%���R~���
�;7�=�w�bj=��z��ؕ3͈_������7���溼Mm:[[�o<�#�������Q,����5�>2$��d��d�,�ʋ�ya ��Z٧qx�0�5�_8Ss_X�j�����2;��)�;�\�h���\f$��
� ?��=
�s1d�jv^+�w9��nx���B(%������Мˇ�Qq��n0�ç�
��r�˹)7��ݺ��=�Kv�̺���������=$��g������~�d��b��A	��8�U;q�&�k@��6���0�
����: �#��S��{��fs����uW�����sh]˶.�T�4C��|���0��X��$O���5���.��U�rM�e�؞<;�}���	,MT/��E�}�ml3�nRS�$K�P^�3���v�V�+p���|��u���X��@�̴��M������^IL"Ĺ�n �F�7	���2�g�}�������_[��J:&��Ml#�.�㿬�B�}�g?�u��Ѳ^�����"�l��6��������"=�s����Eu�=E�����tB����!V�6�_������W��r��+�{6�@
��:z�1v-I��|�Ŧ�E.�ҘT��cs��K]�
ںó?Jy�=WӡN��(�G�g���f+��� �m}�zV��+�5�]�
6芍����UxC�+�6`��2�3ý��L<+��A.?�CD]^�|��Xe��5C� �}�*i����vK+��od�q���L���X�87(�~��[V�.�˅�T�o����+a76�[ǝ����g;f����
n�����m.�z��|��k�'Q�l�	|Z��H,�344d��`��6|�8r�DFi��	(������k���+4�C>�$.����Q"<���[�
7��9� (�Vj�J���Z5�a>�Lzc���
P���ȡa��6i��L�a?�
�cJX�s6� ?^tG�
�=%��ч�9'?���/Nl']a���W�)�*��r�[|��1��j0@�C3��lgz`+7�	b}�v�5���w9�bg��׮ED�_0�}a��o˛��\���F�4�¿S���@��>�k��A��/��$���27Z3�K�P��em[����Y3�E��4qj�_Xb������5OIM\q��D ^�x��d�����9��������=�M���1N�(W"?P��B�v�
��\��"a8�;Y��th��q��|��q,x���M�?��,.���:��ny�;ҙ��i��%���V]��֮���
Ǔ[����s��ԝ�C�~Q�5e��������~�ID?"s�`��!�f,bF��d�7����R�M	�=� r B���I��FVSv|x���4#1�'mO��S\��C���@�ɣ�t�������g�#,�A���kɷ⵩���)��!ۣWfD|
W�v��_���nd�HD���BeR��p�}24�N����}ۘ/�EXU��ʲa(����\5{$S���-Q��W��c�ݞu��M�� �*'�9�?	�[Ӵ([b�FHY�'�x�ȿ��jȨG���:b2���3�;U޴)n�A���+K65��?�l�`H��$�h�FN��������pJ���<Y�>��G(�j�JKs���L1c}���{w�Y�X��i�U���Zs�.�fd��n�񋤛KE�3�>0��������mO� �-J\	�"s�e�2�D�1�'zĆb~�����U���DԮ89�6$$H�P�b��L�*���S1��~��אqC���ָ��9�u�<�v��9G��V0Ϧ�l����M�Q�:"K�Im�/O �.@0��%�5�J�c�I���P��r���P.+2�Dqr�ѐ5C���D�w���q�m�;k�
�=�꓄Y!����I��wC�ݏ�҂����l���>�/j��JY��}`�;�.��t��{F|ޚ:����8r�(D�i8j+Yp�
�aj��d�g�̲�� �6�c�t.��j6��A�Gό�2����4[F��EW<��$�TVWkgQx|�t<�%XF���&��9�x`"���u?�{�᨟��u�D�U��7�^���U�ᆪO#�S�k#e6Ikq7�z�ޤ6-�i��1�0��1q���ts�=t��(n|�8>x�0E�|~�6ٖĸ̠s������ ��L
�R�[�]͉�DL��g�x����5FL1�<���[����ɵ���a�=��ڄ��qM�r�',��2�&i3�DB��L�J��=J'Y_\�� ��F[MvBx*U�>��������W^�;��>x̰�T� H�VW��Y+�mf�r�@�t� ��/!�Y:Al�U��J&��{]�������),cL�R������5܍zv�2	Il�h������80��s��!؍"��@�`�W�����T��'��za �,�/�9�vU�{_�KD�۟?%�h9ԯ���ͮ�n3��|(Z��4�ɶ-{{�?�xl�M�5�&C}�� ���{�[�QL���C����'�����iWc�3�L�n�*��*����Ί_��&�b6�9x���2�r�̭�m)���sUYk�����.\SI"��:Z8`֐��� Y�j�]0> �	��=@�_��t�z^�R��v���mY���?�Ԧy0����I�[��,�U>��n�ǒ"5���D��L6�m7�X+�%i���K�"�ץ%-Y���l�w�����ǩ>H���c�����u6��zC`/k
��C���۾���[񼍑>��W䏜m ���F:*���"ѐ��ҩ�_�ݪ)Ly�T��+�����K�E��d�[>H2^	e*u��_記��N!�0�+`��
*0K�� ���w"��jo���U���綜E��/��b�J(h�.�U�ת�G �~�]jQ�H��9�	M�f�'K=(qoKZ�4�L`/��aU��Ƒb�QJ~[*h�mE��M퉂��ퟞT�E��٨Țf����@+A�I����a�N�hs��]��W��_�s����֥���N�����w��dsɧN��Ô���iKr�Z�;��L���r`�hDgY�C��\�l��q=��qc�4�����'@҆Mq�dm˭�ۤUk�%'O��(l_K���w���'��YO�-���W��]cU\V]�<����զĐ�8�؞\�͜�0��Y#w���P���ې�;z��I��nV�O��2a `�d�vJI��݌o�k7��$m��Ւ�0�$f�A�^(�IS���Q��P���(��顓[K���}�������.w_K�G+��=���*���"��wR�"�u"G�[Y�o��1rHDك��9�Ԏl�L�&�M�U:Q�`�"c�W�	��~�b��j�i�p�C�d�'�B2��Q}(A�u�kU �NK���w򈭌�b$��6�K��"�b��9��)�k�9m��i���V)�e���E�=.�Aׇ�>ˑ�7�Ő8ٵ��l�g���Mk'�*�xO}�a(���et������x:�`�9YR��� �7�g�"&��&�Ad��@l����H��H|Q ��,�/
^@�	 m�a{�I�"v�\�)�@ĐWR!�X