XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�e�}���!��,!?���o���j���%^������!�����j�p_��*����4z��?�S\�H�DW��� ��~]+P�����Z��=�dM$	7���2F5i
���:���&��AR")�98�Cs�Y���!/�UP%KYk�P�GH�h����|Y�7�]�o_i���VC�Rr�T�3z�7����J���Â]�KZ�<��E�p��a�/�=I.XlE[��F�o	uj%}��>�}�xNDw�*�)��	G��4DRWo�Pv��"11+4����K������2��������h���$7C���ɂ;;'[^D[u}f��8�����&S~�r�+�At�Iw�(�ܚmD�c\
<ʑr���H���B.Su�I¹d�L�n�s�����mH"c�UY�J��:�:Q\�x5�+�&g� �G?��Y)�Hƴ�s%��u�0�[�tK�!�A�F�x��L<���<}(+��Y*��M�c<��<�
j��~v�+�<��p`��a��Ǘ#M�}��Э#���9��dQ�����X A_s�SV+ed��
W���&�L� D�%�?�����$���0�aTIK��H�����@����TZ	t��M?���?ፀp��L�'�l+{(�u�+/�ʍ����:��_<�e������{(�iYc&�6���D�������|�D^Wl�8+v;z�>x��1�^~��~�H��l�v3	����]�
���(C��x��z|��<�XlxVHYEB    3da6     fb0t�L~�k#iG��_|3������jro"���p�D�M��Q��+m(�3�2�
nN��jR�N�%��>�o�����ZrC�p���a��qց7�v	~����)OǛZ��0a���yڭ����K�M8`��ZI	��]��B�$]��% ��d=8~�eޠc��ɧ)Q�D�?��+����2> �px�~��K"��ԹQ2����S�p��NG[Ӟ������S�򂋃
�r�����s������c��v���P"�"���cݫ9���h�r� "|}ۤ�~}�ڄ�vΙ����B""WQ-#���q#�gݢ2e�7�~�����׫�:�51A�r:X��sQZ#�?�>��P����a�I��Ey݄�TɎ!�e�QJ�'Z3(�Э���
�"h��a��\)��5Y��+
��j��-Օ8{�%Č��OM��ˌ������s1��YK��.��k_��2�ߐJ�߀>j�1�L������S���ea��GV�f�{C,��z��H�.W�J��oǥ�7��2Gm�C�y��	��{�S�A@���tC�J��u��k���D!�>��"5�kv
'M���ͬ�_���������0Wu=|)o���W���3M/�28�+;+���SZ�w���lӺF@���Aj@��m�c�@l$���ZF�e��ӌ^5�K�Q�$�]��g�i�=�ɖ�Ċ�Qr��,����Ƴ��.��_IvY�4�l�?�l�7�Y�{�-�W�^���O
��=\�S���^ǖ6(��j��_�!D.�T�N��b7��,#���*7�xa��Om�6~���%H3cr��|k2������J�aB�'�6�DH��'�gI�..P�%����f4]c�=�\��[W�\X������t95�E('�P����hɤ��tn8���}ۇ1�CA�r� E�%���*���i?�_�#:'��-0A�=�1)�c�ɯ�#w�Ņ+�e�rn5�ӆ��V�M�Pr�'��^WU]�~�z��P�&W0���`ں��|댏a���'�U��
�������t�\sy���3��x��t�L���$��g��ِ�@z�����jԩ��o��դ����riܝ���|p&�pO}_��y��j�da�x,ضK��W��`�sI��gqpk�c�X�=<�B���>� 0_6�L�����	���mˣ�9>��51`9�?H�>>�#z��� ��3��e��l�q!$�8�J��������(���]M{D�� pyP�*��pꍏ�|9���]��2u>���>�!5'(*�ux
�N��V��^����� 0x�Ff�5Y��aCrK����/�݇_C���<�,Jt�t�s�c咟���u/���>��!ب0��R#�@��']as⳻P�UZ���ac�7��İ`5RF�����@�<'�8嫑r����IA/a�^��$�n����&�/�7����u	�:�����j{�����C�:#6�+���3���([6��^_k�)�zP��Z8ҟ�6���N���d�r~*1��ʶ	&y$��Q� 5�����3c�1(�3��f|?iHz�mF�yb��U$�%LD-��Gx�o�a/�)�8�v�|�[b��(�Γ�E����}F��C���|���9ze��N�EӮ�H��

�g4_B0x�@�Zg���'�g=��.�ﱌ !����[ �jg~(���>��f��h�
��u��$��J�[N=c^� �g��&�1""�	1X�IQ7�A��x�q9w�Z .��D�$����b=Z�8X�L��Y����� /��|#�w��QQ�M�VV��X`��rcl7��8�
K 3l���~�N��gF�r��� ����<��[�"Npl�&+�ܼ���\șE��uȱ��ׄ��bk��B�׼�^���2��+��̾P�т���v�Ψm���L�S�Ю1r�^а��<&�E����E�����1�`���*�� (ϨX��ؒ<0�(��W6�Ԧ"�s������H��R2������M	�1a[,^��L+�H{�$n����-����~:dxN��s�:�wZ9���0.@$\�r�H�����^=���(��Đ��$`dc�t��iJ��4�IW���n,���T!����3cQf���I�zkN�S��悥�N����Lt�Yx����j �����,�&�Ԕ�.Y%�@M��d@��P��\=�Êw�c: ;����B�����]6L�Y�tbd�������������(�y��B���h�T2�\U�����xa���y�n�]iq�V)�h]���� S�0�4�O*� E���'� Q
6y�0�܇G�"%���w��zo���X§P������M���Y4]]�2ժp��9F��h�k�R�J -�D7�)H��˲Sixm�S��_�u1H��r�|�K,̟҈ք>�������|�����j%U�ā"S�t�;���h���[���7!���
���Sa��0�m�d=���?��8'�<&O��k��>Rt��Z�Yk�9U6�B��;qn�P�=�̤[��1�Z=�Tf�sH�)(�����Fu���v%S�Z�|��.b���ˎ�e+��LQ{W�Wx�\�/�s��@c��|�Ʒ}�0���c��|�M)��������_/��6����Lb�)x �J�@0��搽�/�7m��/���Ki�]$yVy��O�X�D���|�~c⅔]?�|Ț�u�3�J!�h����q��M1��nj/�W��B�T9D1yb��ΕjKK�9^-�AM��	�P���f�pٔ�i���h�����K6�f���$�O��,���~ס�bU��$�&�$f��,��^��-yX|N"��7BN�\�>H-U����*�|��h��$%����K�����l����Q�*��o{�
2�X�]��x	�p�B�D-T�r5H�6���hxy�&���ؚ���z�+"�|Yl7UG �?o��c���^��؅�
W�iy��0�"~�+0s��t��S�[��
a�p�]رt�K8v�� �߀�M�rW��v̎]tf��Jؙ"`���A�c�v8�Ϧ��Y&��^�{�	���
��l,�Iw�������bo�Ί�|-�>�"���~J���y�[�Y��Z�к��q�α�kfK�Ύ9#K>3������c��kp���A\�ߵ�J���ݰ�ȽY�[�����QOw��<�a�8sA�7�Œ���+:�i0�.�P���M�s�}j�dj��]B]ojy����jtyQ�-�lIp��j���9���u��)R׻�D���yQ�H��Z1ʷ�Ժٟ�3E_�gS�!������B���F���":4��;Y *�[�+p�E�/���+���З��f�)v��j',�/�
�m��jd�g�x�,�HQ�7"ƽX�CY��G�<������#�p{�(^�h����lw�!��`7�����r�o�	U�{8���~����p�h�e�@,�p�\2��fg!.�,z����� �
#�ai�I&��'
����e����ns#V���vdW^��}Q�I�(M�Z�rn	Sy���RՎ�0���H,����v�R�é��D�d"� AY�R��ݰ�hئ�k�Ȕi��;	@�-/AP��?�P�MA���(�oc�HnE�o���J�(��,=Kc�<���O ����n.{�̟Eb���e.Ft@�6�L��=��b1W�;��U���@�=��V�!6+�h���©{�s�����H�)2�`="��kA�Զ�NL��D�"���T�� ���F���>M�����ur�m������2;��F��k���N�X�Q���&���m���2�����9�A�Y��fH0ȇ�