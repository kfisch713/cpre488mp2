XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.����q�I�����t�3t����x��/�KЊ����q��k���b6�wQ���>v��v�\֓��9?E�Jwxe�riy21�ݵ�����/����Tw���� �3r���#���w� :�(����߀J�X���<7�@d�	
J.�@봎^���ra���+�6�����,��#OZ�%���7Їc��[���9H��sR8��C�Z| -5�c_��%?�Z��gQ'�N͢��� >�.ѧ)��L�C����4XZ�n���@�ő�O|�>0�.z��23����`�����hNuh�0͸�C�]7�3����h��y=ە��� 򐱶�zj*�-8W�@\�NnY)�{+�P��ln9PE{��e���_i�ڗˀeL��fL��h�1M�#mM��%�~~�3 H�*�A_�a�ݤ�n�V��B�aJvD5�:0�(T������n�ٚm	��Fk5+���Uk������mƭ'�^��,�!�d�lm�%��O�t����5��k��F"���_�
_�Ta�e²Y2I�y�/�J�5��1���6��>��.�* C�����e8����3�3���C�@��+
�;�ӱ��F��Ŵ�l�bs�FRz��E2d� ��!��p:�(�j&T9-��G���3U����⫆E�T�qn~�+z�݋���mr���XQm<����m��=RނRL����0�t�N��(�ql���D�~g�it�<vg�vH���XlxVHYEB    893b    1e30~���[*.V��2�v2�R<��b�J��#ͳ��k5�S��Ţ>�bF7��	��u��ë�7p��t^΁�Uߙ|ʏ8��ؕ^�Ú	�%C�����=RI�y"�R+�n����	��m�פ�I���:Q5�45�Nt�W7�  ���^j�F>�7��%S�Lj�_�j�yΌp�
�
���r��<m$�k��Kh���#J��sQwu#��W.;������1�ZѪ�l@bɘ%o���:��+v���g0-z�IaeM�#�i?5>I��V����z�Pa�l.���,Q����7c�D�I�/�8�C�ˣS��Ip���f��)^�'�u��~{s���:uVSv��#;�t�fTKC0�
��u��o����%.@�V�b��S_|�失�s�D��c�-~��
e��� s��&�A L�������-,�@�(��M}7���瞄Y<�@gpb(w�{� W��wAx����pA�?('a�Q��tcJ�,xxX���m����T�@�:��WF՝N��iS�����Mw@yk�7��%�G1�+������_FpЫ�Mk	¢,;������v(�?�m��!��L���/ܪ�����`�>����٧�C�� I��uf<Ft�tuD�"�D�7a�.�]Qn!28QVR��3}<3�~��=�r�Jgì��n��q>��b���C��"��K���hT�5��:5t�*���s'p���	0��@��BH���z��������b&�zX�����r���+h�ȄuU�#�m�������莙M�Љ�E��a��h�XPȱ?V�2=*\���N�ń�XR{���%�Յ�cͨv�x�'�5�Hp�!מ-Z)e遺|J�U������(�E���B�4Zt��Y��Ҽ1{��n��J|��BpoCS:o�b����jK�	���y['�9�-������l���� S�堾�.ϥ�wD��~�e���%��Q0���1�N�WX� 4J�&�M~�,��w�������?'Y��r(�;*A
O�d�:g�!�s������d�r����7@H�->=x�DS�D��{�tꃸ͙IlP�۰i�������4�-�I��J��G��;	xaC�L��V	��%/\�2��l�mE~��H�ъ���_-ZYpK��>(�4�:lj��{.��)�|��BsP�%_&h˫�{�א�1�V��B��d=�1z�K�N�B<ǉ�a�vi�-�
ᓵ�E�sݜ'G�/�O�y׸Y���U��L�:�����!R��<Y�@��<�gsF�uG �:�8�_�g��:tN9X('�T� -V�SHUG��V/v�n�D��w��i�z�9]����/��/(r�-�L���������G��=�������s%��7��XL�v%�����U�k�@���޶�������G�o<��S�9<Ri= �A����Ϛ�KB�qS��Z�0�C��{FyfYQo�h:P|	^���A�on����x oݲ��u}.�Pyk���q<|�gv���m�[B��&�����B"�L��|U5Zp��4�"ۼ?�Zx^�^��� l#��򊳰oZ9����m,V��XD"������8F"��H�:�t�c)�fG\��S���}D�4���&�RxO�g�r�����Y��O��u�����)X��'�fƻh� ������"H�8>U�^�g�;S�>U���kK�r�J�}#�%���ʋ��'=���,����\��"nB�HѐO�m�>2sܔ���߈�P$?I�hy}!���2���ׯ�-���׮����R���1�gB���J2\�K��x�ˬq)��F#8�
�%@��Xk�ؓ��4B��`�wMTp�-r?X���3x���6�U�p����.X}Q�.���GrS�O�5{��SgN9�"���Z={��j�U}�P����c��5iҬq��7]�kz:1�Z�#Nt���ƭFn��z�ab#U ������|vG|�zm$O2�sѺ�ƀ2T�-14�o�\��Ǧ��,�
��Od/Y53}�)Ee�cƿ�K?�7���"�zwe�۞>ߚ�T����+#��ҁ���7�'G�`���AU�]G�=�8;g�O�@�=�{���l{�G��. ��?���Ҝ	;8rh7^�`%��*�B\�����3t �F���z�R2	i�[ؒ}؂��ڜ����4��5Q���"��j�ԣ׹G׬�v[@� =����ԡҨ��*DR��z��=3aX[w�x��{~��sH<O��3��lʎU�Е�5T������p;(s�¨����7<�����W��Ėn���a+;��_W�n�oV�8�ܝu��Ǣ5eA��촉�ۜҿ(M,3�cl�����u,l��qL"�P�5,�y���A5���\��ۮ�Bq��OI��e��.J@��g!�Yƨt����7��P�
�v�)ߙ��w�).�{KQ"j&��>
��a�:ϩVu��Eܣ+�(���I�e=u{1i,8*.	(J@z�ݭ.ǍW�n�A����x	��Z�eu؅T5IY�-������:~�����1������Lj~�K�G~���p����W�-X�V��-h3��m��E��������Г�H���h�E5�x)Fy8��+����@���X�恬в�G���|U|Dd�Z�����Z�O����dC���Q$f�`e���X, uq&�k�����P)H%��PNP��o�⪩Z!��wN�U����6�ƑB���f]h��PZ[�ru�I�s�9���A��E�q�b��Hׄ���7���dxܿC���I������~tJ'�>Rz�@����g��^4�i竾�[{BY��o4��A�?ݜ���[�T��@�[�|�q"ʃ�]����8RFXK{�H�*�����-����]8�(E�ns����A�9����z9\v���V���OW��H�m�s���T2H����P��Q�wS�>��l$Ld������s�M�օ�F�{ô�Lo՞n��.���oΊ�د���4�2r_B1��Ap�^W�oz�B���sH�f<M������ӆ}��GA~�Qps&�n����5�@p��m�&����6�Ү��\���M���DcI1�ҫ&���@ꑷy��z+� �IȀu��ADcz��ά��B_�4��R`���3�G��۰B�x2y}���ZMH����yJ�?&wcZ��ʝ��Z�m��~L�RZ�:Ծ���ޯ�|�D��H��;�R�(�2?o�Ӭ��r 8�Qv�E0�ͱl֦Bt�#���`��+�L��Nj5��l������]��&{����}��i��0F<f�+�B�p@���!j�q�%"�������mX{�1��Q��h�N��Q+l*�Xd�a]��ʃQVx`�����O��G�@;�AWJ�G,�O�q�������d@��bkI$��l�O�H։�2�Ť+iF�YўLh�u>D��@���V��.���050���ލ�,HX�O+ܩ`#�^ �8yQ��d�&?F�S����7/'����ɻ����6	K�<%��]�����}o޴A�2�3	pZ�ͫ�n~-��zq�\��%�+1���u���3�-�j?�������Ce`ᎏ,G��
wت�3�`�ڮ�8�<w�r�J	�F98i3j��gRԯ���"+�2F
���&����.��YsZ�+�_��U��^����	��zL�e�N˜^��ן�kS���QԿC�{��fRgo�`y)5*�@�H�����o,�8+a��!��1�}�{iXQO�-Yx���@Jy?v{���^	�ňܓ�]���N5��rˁ�77-h�z�
�=��m(��~a�w��V���������ۘ�JC�W�*-����b�k1�P��1�y��&X�G��<!���N��+��z�H��M"����~t���/☽߬�~~����֕��7�l�����+�AT�HIq�W�l�$* �Y� �{��RI+����.�W�bx�$��88�4jyK� ڭ�]PK��آl6�P��O���<��;5�4�|�ܧ�䕢�Z�^g�9 M.�p��L1�ۗ�Ns�_�j��<[���T=��$C�ܰ}yl��/�Vƭè�~tp���G�x�El`Ӡ�����}m��D��{�<���e�����S�s��7�M����~�R.�W��~g��HOb���2�X�j��Q>��>b��ѝ�C}aW�/y��PQ�@���������9���S=�e��飧��Ks%��(x�]���ɔF��~���s��D������D�SBM+U/+(OOz���ɣ󙻫��۟�4�4���]��Axz���u�G҉9�@�h�>��i16Sʒ.{{ɉr͊����V�I�P���0ϫ.��ے��Z&j��(���ױ��`��+�V�8�r*�FΥ��`V�Zꁉ�/�pN&��l��n4$@�u��R����u-�:#�h����W�]�~�vB��sMLK�f�ޔ$0;�K:s(q��sAN��aMt�C!��]5�爛(0�e�Bs�HF���[�ҟ5)�/Mg���@���#k㊨�[<,�3��&ZJ.*z�S��2*�y�5�Q�}u����ރAŕ�Q�h���E�����b��zxO��h�g1f�3H���o5���Ep�qny�X��
��W�q(R���hH��͇9��BF�,�� O�M]S#,����������*���Xb�}n�(������)��a�Bje\�t ;TՏ8 K=Bx��'Y+����	�z�Q����l��n(�杭���Z$!JH��%�t؝���2X�h�Vޚ��Ҡ�氕?�l`w��@Ω�Ễ)M���?~�N�4 �ʒ�����.C-�H��E�5�@��l��2��r���7II�����I���~I�z"������t�\�[@�я���a���;G�N(�%�x\t�oܤ��>T����冽NxkjZo�\9�ݕV�R	7g"vzB�Q�%y�K��Our������Y������ꊩ)��R�T�B&�L��K��ܫ�)�2ƽe���՚}�O�+Ǻ���\Z�u��������j��3P�����,��D3ɿ�^�H��/�l�.0.LdVC^��sg�XΝ�+r����''� ���Ǭ������R��8���̜�$������x�v�P��j��]��H�J������BEF3�)�>�N����R�mሣ�q�Ad0�q#���m���!����*'�
��=Fʫ�\b�^k��J]	�6�=ٷ��cnZͩcda���t��{t-Wj���ɯ諭ۿ�Y~���Gx g�>����߭ �ZT�\���SZ̖��-Cz-���C�m*�D�M�����*�e���cL��[F�AimIK`�6���]2�^x�>��&SI����̃;ls��ز�5�����$�r�%��o��
�r��	�b�����IC�o?�N�Z02�K�����i��d�h@�t$�h���e1����ƗS���Oq��NeE;ǀ@��t�a�s�y�X�l'��2=�����@�y\6��ב����7�bU�,>�Cɶ� �_�p���U���5��\>>�B�쭤?<d��T�$.�>������a���x�����7�d;���l�x�:�����]���I�@Zڏ�sdjU�(ΗP�\�V��bUL�p��c��n�R�K��]
Y�P�yӹI嵟O#��׼"3�����3�	>�v��0��P �2La`��3�0�*{���)��8�s���{�ŝ9n�+5�g\"�5��Qޔ�쉕�$����ǻG��jÓZ4� G!�Eh��=3y��i���Ojs�:]{��(�)���Z��L��!���(Z�#�G#��{Q�ř��gk�^�u
��1� `ͺ� ���=�.=�+4#0���UH�n�<�Gk��n�cJ+�~��tz�sE�@^�P�F��"Z�<�	�&OSɐ46�&�Dn�*��R1.�/(	�I�X��dAz�@��ff������ɝc95���&&���褕#z(��U��uP-�;��L���ۢ0R-�2U�r���5 .�������#���TD����y؟��We�t����"���P�����aY��|֫�oLX��3���:��Oy�Z�nz���LP�(�2�aɄ0�_#�)�U��\���o4oQ�H.(�Yr;�n��fI^@�"޾ijS�(Ba����Cj�J���!;�rU����
�8��-�:x�Κ�r ��lv��L�.��L���_�_�^LZ"���Y~�K�nG34�wUz���^l���sWB��ݣ�'xr��sn�X����bI5�z�E�m�+3"rJPb�א(�".>��ٕ��3�z��f�͹K�ffO379��N���|�b��d�q�oj ��x�2�Lǟ�d���ގ���<�h�P.J��ZH�T���-�#��'�CU3lo�o$���Yʄ�pV�Ւֳ6ON�>�	��w�_�V�rI��4���%�h-��x]��X�a�f�֥��`���Ј@�v����C��������O�v��������"�y�������0pƍ�ۿ $N�M�����~Q��a�� �=���c��.����mٕq�� ����9�6n�t�̐�Mȼ�����F��q�Ap�E��ۢ:~"X��7j��﻽�[�g"�^U��+qϚLUoY��@['�XFKf��H���޾��68�^���6����XW���l�Im5%�?�p����������1��0p�uY2�ÀX�'�ꢏ����^?2@	Zcΰ��b�oF�1/`cG��_հW��h���R�����V��+j^Kz�X@���-�X�Tp1Xx�G����e�����h&A�E̿=��iY�?#�gu�L��
�7:dA:�Kp��G�9�r���Tg�km�s(#�
��a���6� �>��ym�6S]��	2�3k���:�̠� #z0*,�p�����٩Q��4f�kf��Kl!(��$F�����֯<����0��km7�.g���f��)$u���ͥh�ө�~ذ���$
X��a�i�k�<�8&��!R�hRPR�"ZY��&c���q�5dM�͗�!Ң��$�v<��u:0�J�K%��EC�열�vƤ�8��lK�@<c�=�ږo���&�T> a V��ÖDvj,(�]/L>/*���X�y�:P�t�B�n�B��
�ayl/	�O�1���K�EF����>h�wM�RoCX���uAg�b�)���#X��
n�p���R<'c�8��tY�i�ӌ�
�`��M�g-B�����[�.��b�㳪F����D�*��;	Y%����2��ܦ-��d[��Ԡ�䃾AV���4��a���ì���ٗt�<f����>A�C�)6�8�N&�x�f��2
8����kz�����C4�a&S�F���{���KY�G�=n� .n�b����#�����?�k�i�<�x7�+�o~�*p��z��W�gs��s��jg1��M���I��|�f�^�"Ӿ2d