XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���1��k��m���A���#4!�B[-�]�p#	���g�릂ϝ��[���1�
l;��a	Q4�N	��JJ� ���y1_�6�-P}���X-l�CJd�ayF��I`�A,q�^�唘����k�Ӊ�϶���*U ��v�D�0���u��1�����+�2��bz�nW4hI�PK��N�ӌ�sC�Y-�¡2���f��h^7�mC@� <��l���]�ȍ�!�l,���r�CN!������4_��jg�)�,K��/;ǘ��;�j����_8�:�h̨��Ό���+V��d6ʞ)Co��00�g�e~|ˈ�u4����rp� �l��:��	��u����7��KǤI����|�GEp���֫�e�~sN�s���ZCA�����Y�o�[C���5s���*'���;	�#�����������U�5�jޭ�)n�;6HS�Z�P�3Z�f��{~H���_�,�<�/D��&k5DlL�0v���%醀Ѷ��238؜ZU�����������I��f��\��H���2�|��~?���ǩu��+��Q+�!$-�g<mU3���=F�{#�����	W��n�3�Gx�tsΙ���u�� ���!J1-몼s�)�F&RЎ�Ќ_�=q�k^-d��u�ͧ��Op�����8�T�[������ØaҠ>�X?����UlY��uZ4,�5}��v~�F��
�n����Jo{u!VI�R/Bo��nb��n/XlxVHYEB    3e93    10b0U�7f�|.�@ٔ���{������%�nAƨ�e뻛��W�M���#�_G��	l(�/�gnP8@��I(��:U�M5�[m�����	��bv�:��5[�X������WW�<�hF�G�S�+��K��9��8� B<{��.�
�e��\���\L� �7iڤ�������/ޖ*�a��'�Q;N��J|��\j�<65R:��H��/������Pu�R?��5� ���"E��� �DI���ü'����u���~b$e��p�"�;��\�žWeu��v��J]�7O�)��Zg��hZK��f3>ǫ��H��f0�?V��i�өR�JG�Z�S�hKJ���oQbæ����<F��������#��8��J��1R�T| �
�7aL`�
�&�@���L^����dGo[�8	����/U�̀�_(�7��#L�8�X&��ޘ��ѿo����I7VDr����#Q�6xp��V����Wt�@�Vr��߾���	�V�
���"�$H_��[�0`�뇟�@v�=�x��ZU=}�稉9>��MЗ&?���Y�{�����*��b,�[��i`Tz�B�{��֭����w�������hm~Q��+�T.'�Z��F���@ٌ�t����YSV����_�2�Pj]�=�*��xћ-��҄�(Z'�.�.U_2b��Eb���T��H�/�Ѓ��jlGX^�.rc�<���x�W2�Q�+W��9�QC�=S͕�|i���o���4�QS�6��R�r�)���"�{9�I�\���H��m��ɊȀ�9.�whK�����Cl��r�d؆5i
�
2o�����_�p�72�Yrج��0Q:�s��}a�����D	!��bw��C��ԝL�Ff�nu���L��	��/Q�*��f�	ZtZ"��!�q��;��۽��z��S���KwÂ�U+��I-�%x>+s��U���Ӥv�)��.r�ϟQÿ�@-�Z�J��Q���������;ӾV��8�$`��(�`�DI�|�`�����t�4��w�$Do#mր�L����o��֍����F/��znW3K��{�}��Q	_v�
�7�����z�D��2�!�G$�u��_Y��uu�L/JD���Z���_�U�?»�. �G���	����{��C@Z�#�6S��U�t��m �%�FG#�i�U�V*i�W�X���mS�t3(f��w�wy�+����m��j��:n��~Hd��S#��4�����;Lɻ�f8#7\�|�2P�y��K����Ke��m�s���_��q-��4�#���4�����1*�Ѫ/I{�eQ3~%�9� 0mF7�[����_�|b���l��I�D9Uu�<LՍ��׺�M����sQ
U���K�I��<0Q��mE A�<��W
w˩��'��<pL��JN��:��M9[p���>�]u�U��ZEZEI�\� �h��)K7�ة���a�4F��F'e�Ȋ��^�t6�h��r����	�����,2	�i��r�"�M#� ���e0[G������\h�3U,x����Hvr��@��$�aiȖ>y��Ry]}@���Ē/2VY�Q��|�3�_:^�/Ц�����#��d�%���ʱ\�eU��_f*V�,�j}0|�#֦��5QZC�7?� ��؉�W�{�'�Ӱ�K�u��P�)����%lG��V���&�\�y�ާ�Z�"�95�EWc��qGS������P0'���^͹���c8�D�@b�݄������~� "r���y5��v �w)����Z^�r+}!o�q5o9A�ۗ��Й_cJ�P7��@&�#���/xy���)xϽwOm.�5��AU��@C&x��{��i�(|a{�n���~����b�ާ��v;�#O,�ϯ\)qBc��⾅��!����$q̈́��r^|{M�F2�h��'��`O(e\7����PS�Q�i�̸P��YOݮ0SD����D`|!\����Y�-�PD�p�;�������>����Ыz4(�� 4$�8^@ �r)�p�}�1��R3։R��K̀�V���j��9��?�8kO������.�aS�ս�r��p��y�Ӧ��(�kpH��Y�_�L��m��3��x;���}푫c��y௫��9&�C�k�t�:CR�5�_6��q����������ŏ�����^
nڗZȵM�cI��+N�~�{�0���/�ĥ�'hG�N�P�mF�D:K!��u���RHE��p�kz68�m���_��	x��SH��V���� ґ��5�{�%:GGt�1�7@4�Ɂ�R�0��V��{ڔL�t�i���������Ϙ�RE+�=�d���Ǿ�+�u���������M>��*.�L=�BQ��drH%uLVp'@aɧ����-f~3��A�9(���v|x�t]��h>�¶2n�ҽ9v���\�d��¬^e�*�A�z[���ĦQ2�n$����>~�|�\�Sc���?k�DJ_Q08��$��e�d%~}~v�;�}�%�n��[x�˕�|��M��Ѩ�`��'iC��+n�]������-ܹZ^Qk���q���ae]�Y!)��~��2���%�>��g�����t�������TAyacp�%S6��Hz$�8�Bڔ�������S9(B���g��-gwδ҈Y=S*��~H����6��� �����[|�ʸÌk�-���2��O?���՜�UٱE,Ҁ�'�������E.-�S8k�Ʃ974>�,���JIC_�f�Jj���HVcFlFb[��=� �N`g[��m�*�7�K��� rM����%k��U��Z�v!Ԉ.A�>�H��������-L�>�d�+�ֵps�٥,�Z�����3oD�Ę�l�/P7�ZmA��hF�Z��֌Y��6��l��b�Q7�u��aɖ�՚�MXM_��$sr�벦�����1?�+%���8��/�	����9<�n���K.�_����G�my�GT*�Z�-SQ�:���~S�������.BZ`�p��(Q?Q����V�#yL��+;5�k����U;U��g�GTr;�WꞇC���7��v�y��N�^�����s�>���N+Q��o�3q��H6%����fn����|%����ihYU�����EX�IQ�sfӡ�볨�߁w���ξ��>O����8��������?�!��¶曈8��� %�G�H��μ�]-CB��T��4�N��&H�?ȸ��^�fÛ�Pmwb5�c��5Kv���;�M��2/f5��d7<�pyB��ǢD��F�$�V�:Q�����)n���O�nw��Gf��?�z�5������ct�T*���z4��(��.��V5j��J[6:��`
��Rwr+��cN��>z\�	�=�P0���<��
h�����U|�F/�_����>'��Bи�i�"׋|�ܙ9�^+��e擬��<�q�GAX�����ѐ2GV���Q���̿��|kGA�6]�9�)E[[��F��Cv.̌�ޜ(�$Qb/ ��C�\�U������N]��^�*��� ���#���LO��1��c�Q@�f�+/3��s�����\��2�@�С�E�I�P��������@���ԵxN}`����Css��g��6,L��WS�W��F��۠��Z�)H�P��r͠�ϫ{��r�YU�r'	_`�֠{��`N-��*q�}\�MS|8Ab�l˻�� Z�Ҳ�t���/b�P#Onu�r!�X�.�	U��;S��%��Y�S��� ����y�Y������f\�vq�U XKs�4TI!�l^�qyp�ϳ�������������tJ�ǲ��2D��o9�\�� 7��q$��E�ڮ�A�ˆ_�bA��S1�z0K{v|&^�k�KT?�Gt$�[����[VH):�p8���Տs3u�pn�px���??��@���w�%�K64�6�q3'vB~�ÿ��m�15�}!�m���oL�R
IkNX�-��G�o�P��9\�l͟�r[K9.�,�ʕO�D�b @�<ɠ��8T�ឿm���H�v��&�u�&����#�̤- P��W_l���B%�I32x����3Y�g�ѥ�J~@L��C1�`$U�%9�c���3]