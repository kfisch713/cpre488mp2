XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$y���H!	�e���{'tg�-x�J���ܑ�'����x����L'g�i�~��Tz����`I6c�� �C�DH�;tkHi�
�d��)������XIUݞ��O�1���(�X8c�D��t`DU�;��vy���'���>േ�A�{�Ҋʞ,����	�КT�sA���(_����l	�x֘r�A=�˟�K�����<kX"Ƚ�������ah��?��Ϋ�d�a���ӄ?I��sbq���W���<F�/,:U�8i��OF}c�����\��{_���I��Oe�VGT��T�31aQ�^_\��j��Lh��ߨ_;��A� ڝ%}s���߻$`R��h�*9�B��$t��6e}p,�8r�eaqڽ�*kJEŀ���K�T[�5�R,uz� �. |� ��砐�����k�H=vƭ3���<c��S�F�Ap�U�7b�)U�
�N��,��9	���C2H��Ik�UW�9C�?(���1Hi�}��l����/��UX��Rt��g�}
d#�P�E=;&�'/��j0h>l��-7�/���X2W�a0}.�޸W ��"^��IS���D��y9KUI�t���\��D�ʖ��wp����,_
ή�W�⫳g�D�f��ޛ[�|������7��*��zf/�Na~�e��]Kj�[�]T3W;H}��7�j���)����S%F�-�y���r�vڠ0U�L����l �&㉤b=��Ћ�8�s�w�U��^�����XlxVHYEB    5224    1740�R���E� ��c�����5�0�>mP'hؠ/��jj5=}V�����z�p
^�7Z����6�bX��>�7�F�_�%�E���x�8|��L�a^Vn7�²����6�+ɶ�} &1r;r� ��k//2��Q����"�������s�DR$}&:�6�l���ߧ�@oi{�J����F[cQ��Q1 �l�@H���+�-?�iv>O��
�ȔF�[:�}$U�/0Q�r����&���ʒ�U�p�&���N8��8�l�-��,�ddf����>��X�*�~<�o֝�UQ��_�q�D�@�u���60�@5�m�|�)�k �IҸ
�;i'��lO�^\e�6u���0!ߟfd#w��İg˴�-E �E��H��"���_��r�u���p���5�CLq��@���,˛��¢֬C��u ���҃�7�K4o@�c#>�&��b�~�U��
$N�vД�h��Rx}��[L�"��u̴z�ô���C:��� ;1�g��|��\����e��w# c�$D7�å����u�>�S����(����PpF�Y��ЀVE�y&:�p:����ժ�PU�X��X^�����[�N��8u���������'�O����(쩭f��$5K�(��>��a}��x�8nV�r"8.�:�|�8AS���av���V���S9bo�Ɔ�`.4ޓl�H�x;��E&�Nר=bHg"㫀L�ۨ�%�?��L�ǅ����3n���z�n�c�������V:�{aɡ��r�>c4�>���k.<Z~��r+)���/�=��X�k5�F-��d"B�D	����N]�	/7����&v�='8�v�m �6�W\�NhX���0�P1s@�^�I�\�J�Dw��ŃrGbɝ��Ml�cd!^Z��"�E6������X��h#aPF$�K��.䋺�R�J�h&��[$4���f\h��\�D�c��Q+�U_�5�-r�z�5��'�c�يg�n��S�@�l�%�፫���-3��/�P��횊�B�p����L���	��,B2�)�=��F�J@~�l�%�m/��kǎ��dB�G*'H�xt`66`��B��m`2���8��%<�I#���8r�_G�Q���f LӪ���4��]5+N�ٟ:�h]Cw�c2-�ՐCG-����ܨ'p[<��xF��D�8��*1�ާ��^9�N>�vH1������u"h�Z��}��z���k����U;͘Ւ7:)I�������Ǣ2�n.�rJ	�4C���w-�� �>�}`E���p#.G��-D����5�٠-��+z���0	�����[�w���@|p3���h|�_��a�D
�4��Gn1��?Z�l�HG�鶋H�|�\/��{v�(��$%���c�a�o�� 8!�'r�o���ZIԅ(�j�=�q˖�#��%��}�ݬ�~S��ߍf̞o�Vz�]�-�}-�ųi�����W���;>�{����F�V�/?�~�"~ud4J*T�?O�6bM�"j����O��6 �N�Әup�GO���j�y2OTz�
W��̆Xuy�x�'dw�ƻ��_G3c�\-����|�T��%O�$�*I;J��t=�"�r?�l.�}�^0֢��>(t���H5�b��4'g��Q,�P�=�Q�5P��-��Ԩo�-6$T���_�ɱ@��Wh���8�q;h��4�6('��"�O:�G0'G��:A�5�Q���_��ʎ�	��$��7����Y^�fh~�c<Q[�41A�cb��.L	U���t<l��DCy]�5G���dMԞt-JZ���v�m��J�E���z�R�Bp���u3���n�ۨ��)�W3�x�Oj�0��0�}b�kb�򮜚P�ҢzPQ���e$�R�������_�ޘ�k���T��o7�Af��=�E���PC?�]N���4�VQ:+��� �V-�dPk�ô<�W�`P
a%���KC�8uY���Q=?����Uo[���h���U���Y"Yo�] #�3Xf�
[y�]L���-ݓLE����.�|H+���*kʱ:ۊ����v�?6�J]S4D[�e�Ols#C��%ï.���?I׽��TxAԔ
L/*�=;���Q���|v��`أ,��(d�e��$mEc��i�)�� >!3�t��9&nF
��I�<�7��^��e��o��
�bV%3�˚�s=�ZB��?�ynw�,�^gC;����М��x#;�A��F� ��iۧ�z��ǽ��}8��u�!��?[�'�E����#��Tx�x�Fꕮg}QU�;�C1{�iؕ�8�)˙�����L�?�pV�H<P;�^mG�I+SP	f0����U;[��Q��삪�W�+m�j�7���}.��w�X6m�=lU��cQJ��}iݥ����w�j����j�U����4�$z��d�y���(!��ϿA\l��J�8l��� }a�AR;l�r�O-k����6<P6G��A+J�N����J���g��@��Lr�I-1��Y������1|(D��>�c:�Uu=B<4U�(E�Ȋr�^�P��B�\��ى+�,pxm}��� ,?fH78`%,�C.�� F��2�u��t�Ŕ�@Qm]�R�1a���8s���#f���Q�
\�rWʼZ�؟F�$�t�&K%�%�C8�e�}E�ƥ3/"o���m1�4?�X��.S��\�
�ԍ��@�<���}�_|�L�Uøm���5,s@y9��J)��el�>c ��s
�7Sq�Q/dSɲ�(-��>V���m%������.���ޝ�v��@B���N��7v56���6��e�1R�8_�<��J�r���`:��Q.�����=}�����^}���b0�tz�^�3�s�:G��;�aI����dst;�<�+s�
-J- Ц���Rsc;�b���K��EO�P�{;�&�2�AJ��=�H2�Q���C���p p�o9��俰�ʞ�6��+��ye�㎌�nI%V�N7�p���p�� v|m�p���W��Mk��Ҋ���o���U���rM��g�t�pm~%��,�����GKnyǸ��--ja��v�h�is�M�/
b�\}���|�����0P2Һ�h����j�Zww=�>�o�/[��>8��%���o�x~�����88x&�șc|u��i\���X5ȼxR�'���oY��O�=�eyp��:�����j���*�,�&S;�J���R<�}t5Z��5�o��-�,\i���#a�Q���	�'��>q�#sn�Wd�$� ˖�z9�y,��~K��Y��%�-� Òz�v����/756>�#X{�(��C���y���4��"�ޠ���S��鐶��m`o������NxQ8���.b�2��j'ꭀ�٠Zx˝��j��*����_�(x� 82���[O:UZ6wJϰfm���K���u(:��[��¹��h����.�F��]
@}^Ѱ����)�
S����Ց��1�\<�@�4����
miz�<L�07k�⹄�ظ�f�Ey�ȉ0h��/��`#�����9�0[�s��m@���I���`x�w����E*m����i�b�Eb���.����:�fS+�F��&�ID��%��~r|PW�K
�=:�/�5��o�}0w���"����K�m����>�μ�c�D@��N���u��:b9Z���	��LQ䕻��T����e��Zr)vOݨ��w�		 8�-�iBE�Kz����S�8��i�R�h8g�'}�7� ��ek��T�&���rZ�SHU�èM����_����>��JH���F:g��A~6��+9�=K�E��Yw�����ܒ��p+�$yj1���^�- 'Q6K�d�6�*<�=w��M����z1�ꍂ:�9N�썬o
�������Npwª������7���� ��Ye�rB���h�-
�0Z�gf�~cس��;.Y��4Ӌ+�|��|�ٸx�������'���s���� �PZ	�(�9S� �z~����1QN�9�}�-��k`P緙Bp��?��E��O\�$"�!v��n�<�#�RtO�X��� ����9C�O#��-�y�f��z'��p�R�j�����m�T,G��꽵eG��>g�[�QB
y�]��������ŏ(v��6"Į9bKW�X�l�ӧ�x�ߘ唽��o8C�+f���	��/���W�-�F��MʷV��������W}=�G��>���Nn5K1� �~^쮩9﬒�N���S7nF"f�S��I�]V�$ȗ}����S��E�bZ:��!���b��=0�d�U���ٝ'eh���1�!���3�E�*�W��88������Z��`t�=[s���i�����ɞ��䐵�E��)�)�iUB��w�M};z���(���kQ�O;j8�S����m�w��'�e��v����	H`�Zfo�O o����-_�v��M_����W�{��;� �������c@�� �X�B���gh�Pb 3�k�ca��qQZ���5m��7_!̃e�|W�^����W8��VC�>�Wfb�́�g��*1��w@��'�K�f��0Y%��5��6ɢ����ڮR���ey"2Nށ�v�[�i"P(�1�H��6��m��QXo{nMmQ���`(�H�b1Z� �Qy�^R��	��Sg�GQ�	0/���[�6�0��:L�ѳ� XL`#�a�<������?g%B�d�}����_�3�Acjt,��Ϧ��͞��A��b����3��5�=g��0$�oB�L�Cn1�)էZ$(駏! G�R[�&���M4�ˤ��OUy��nǺt� �q	��`5 )�#C��S^璮`���	f߅3��-�W�Z���^�g2g�e;A��a��f%ȗ`"�aj#��F�]kz��ڲ��e+�%gPe�3e�0=Q�p����ɉ�U�6��J�3mp��g���j���{�n�M��:��0�"�7�d�I���v���]��cQJ��qʐ�a�ȼ_JF�}�x�6�+c��������'�#+�����r���
'�`䑲l].f&c�(�2��g���e�u�e�ȯ�t��F���X����b���،n�2�`l��Η+�x�V��2 �L�)�	o��g��8���BkN��'Z$G�j*���k�R�D1�)�2�Uq����s-�����[��Eh�(%��O6퉀o��f;��%m�B�q���Ȯ�y(��g;��G�.��.q�7���F�O�Z��{TP֊�
��c�����vyGt�!D쌓��4O��5E���&�R+���x���i�a�8�z�WP��`��.��ű
ꧺ�����{���;K����M��[�?[R��J��Cs)��cg��ם94���}d��m2���L����T��rhޒ�r��f���"��K`k�Z���Ch��={��[mL�bt���+&gFI�ʥHI�%��҇YZ����m�O��.��iT�K��=9�2�(8���d�;ԭ��+`�uߑc�T9.t"�b�ti)gTI���G
�헸�2�=�9a�a��V#�I<���Q��N���4<X/�e�ڍ�sdĸX��|2����IjJX�2-�4?�7	�?��������@� ouJ���n2>e�
�����]�?��u_���Os��Y*��P���:����}����#>=�2nN�k�&y:��ǡ����b�]4|�KKt�T���LyS�\�W��*�_�xE�쑚��2	�U��f|�`�w�ȼC��Gޑ�Ö���c4�=S�Չ;�␄