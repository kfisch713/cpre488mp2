XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-8��u,�s�۠?�l8�%�z/q�	|��ܒW*	�,!##�w ���l��h���ɞ��]��9E\C����cw:�r2 Oe��[�m���<����RW��섆�"����R-�1#�d��+t+g�Ox�@�0�����?XL���V&*C�
`[�����Jk���J�ۘaaw�z��mI9�-FR�6WiCHO����B</�3In� ��I�<���ڬr2�Β��H��l���cE���;�J%����Ϩu˽H�\�GR�U�*<�HơN�ynD�f����]�Kf����d���^h��m�v�WL���i�8�)�|6>�5ݹ�Ͱ��"�h��;���Q�oAם�{�;7�������,O����N��\uo�@ ���������@�����Uէ��4b��\U4��k!�"�Bg�o�����mC��z�M�s��Uy�tc*-ٺ�2�5,>�+���e��y������s��j�� b����|�)�w.u��V� y�����ɕ�gCi�>I��j��E���.�yu|�4�EW�)���B��R=�>�X�:���FN��ǻv��>�%������N�3����9��ߣa;��J��t6�ݣ���o+'G��W�D�H(��=Ϫ���$y7@�x�mc��d6�,�'��@(��#Zُl��2�o�Z�����z?m���W+�@�,�<ŔG���Su�u�s��F�~�Y���}�}9��UB0K�Ş��MHW�D6s1>o�&��^PXlxVHYEB    241a     ad0]�6d��E�I���=� �!wGg�O�w�7min��؉g5C��:)$$��|5x�t�4�����~_�;<wV~C�h����|qv
�$�t]�*-�U�I����g}��Y����i�V%��ɜ�<5oI/�6($�����J}�=��4AҊ���7�9N�ĭnT!V�*�=s֛���8,U�z[kj���G����7rWU��l������&�KPks���p8],�=�T���I'a�m ��� ΢F��+3w��p6>:�#�ڽu�	�޳؏�,%uf��Do�Oz��{Bw$��F���ql>/��ū�=2cW�6��6i�qQ�仦y(ϵ_��{;ѓ,=.�E�;�H��c�}�|$U�ıP�į8����R�����@�0��+����ks�.�<�V�� ;�V�g��s��n��1o�����׷@,�J�jѾ>h#�K�'Kf팾B��	�qe��{ �zCz�s��D��鵽Q�����6Ct���=�u)��l�b_��Л+V��h+�k��W���}$�� �|)#����lޮ�e�+�i�&���26��}��4���������,n���xIO� ��U�FEa9���^ܗ��NG�k��6f��s)�7* ��H����J��5ԟ��֪�hh��h���NIS�/j�&3p�{O�r�

��w�9�l3]��و싃)�(��HU'��
�[�J-��0n�B�B�C��e�U���Zm}��^-�$����/��	o����L�Z�X�e���-����%}���f>�"�?*]���E\
��걬 �����iM���=='w�6ۇӥm{�׵��؋�M�6�K|2P���]��7s:K8~ ����*Ss�H;J=����m����j�Gԕ�n�����c-��\�8�ev���wJ-k���n{�Z5�4�������B-N�Uq��S;K�+�t}Ϣz�
&	����w���g��ͭ�4�o�1iƦ6`\&�`��V;���g�W���A?�)ٺ����CB�%��G�p�j,��4	�CN�i�!n�bvJ����ߑk�9Cp��!^j�N�s�\�q_�/��V4�=��ٝ�~S�`���/�3�v7�ig� \�󙨅��F���&&����,��l@�-Z~�~6m�Hp��-��Hz��j�~��m�$:�AR"�sP�U#0����1Y��e �B��]����Lerh��8S�:��[~Я�P��wz{2Ƕ���`��o��ϼ&M�r�rE1�4�GU$7ߪYC&Ω6���
��&�i1�2�W����-X>��)�������-̢�<a%+�~� 5�;�]�[�=� ���uV(�/Oz�9!��]k�A�z8X��ʍ��1 1�a63�{8��_�S_?\�t��m�J��!6Y�e����̧Z9

����B���d���.�y5lAtC�g�=�cp�����w�iR�R�&�G:��� ��;`5�n�I�z�-���QY\xhc��Ӊ�ܱ�#�5DϜ\� ��.�^mk>��m#.m �O`�o;���NVx�c�[akU:˘���� ��oܑ�c/�)��,V24�(��x���wT���0k���|=�ޙҪ�{���7ǐ\c�V��ٌA��)3.WX��ݪ�,� ��l �%/�v���fB�T�Be=�=�g��.����{��݄33UL)'��7ڵrA��h�Lha��`�����z���,+�)H3L�� ��@�Ʀ�=h��WX�uG�.�ᱣ��C���Q�8����A��n�_��@Ҩ�Me�o7`�G���+�����Q���'�H�45,�<^c��vߧ�Y�30?�p���L{���`۰�hܮ��0(3�YXz�9;����mG\BĜ�,Ȥ�����]@y�w����O�"J�} �F6G��D?�r(�j��D��9���[h��E}j��15�����Ӥ�ox���m�L���X_v��uoʀ�l<�؇��v�M\Dg�$dQ�L]�C�k-�����a����/Ǭ'�2���0Y61�����I�F̞��!Pa٢�c���x'	�$Ab��G)��4�,������Һ
��r�#R!Wf�S� �1:إ-	ͭ�Q[��r�ʀ��W=��h��\���y���Rx�\V4	|ag�HjѦ����6T�fd���s�[�%S��n$ uS#FZ�I#U�z*H�j���{�����Jm�$`*��T�T�Ml+�(7�J)��nf���&�S�hd�}����fXbX�~l��گ� v�;8\���X�-��Z#_F3L�Z�K����\�-�y�٭\��6����36!��UP�V��r���u9a��z��t��^�h�CQ<�T���Ի�g�M����]��%�
'yq[Vk����@��ׅ��
-01�%���r;�u$5�����M1
��g�h�{�s�n{�~���*h��,iL5�����fva������#c�f]����<!-^��sN"=� +9���q�T�(��V���g?b/���W!Ky|p�c
l����T�PX9Y�Ϭ|�%�=�����ɷ<
sR��e���sa�K��^�ܥ8n���h|P]��{��X!�9�R����i��cXk��a�9�.u�NA�@��>���$����Q���F�P�D�yH"s;�V��7�J`j��7���ʸ>���&��v�P���