XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t}��*�6|�}���#�D�n�b�(�Q?�:VnYj� ���oED�My+K�,��E��9wu��Ys�w�F��z�Q�l\�m��o_�k�S��?�Yp�o�A�E𴪘�
���7Z��`�J��9��=���]���Ux��!�x��G2_�5wiu�o��g�!�P�?�Z�x����H�(ngs��+����[����<��}���<R�+J��n �?�Ko���x�Q� ���f�(9��������U���E�Lz�?�l�H�d��|5�F�'�1���W
=J��S!��Ib��B�Tyk���܉�4�b�V�<���S�9B0ƢC%5�8K���O�/WG08UF����j�3�7��F&�S�j1AP䷳�Q-�?��V�!��Z}ί�vW�eɪ�f�e`�
���u�fkX����xηi���# � u�I=Wp}Q�}c!s�upv��:�H�q�F-�{�������x"b���FGr�#_�Rc��z� ��&c�ֳ��)�<j�ז݄��O��@�s�b?#����a`6�\-��������;&�IQ/����/�:]�L?H��ߚ�O^r�+6N0}�3 |�}�D�v�)w6'<:ڏ(�m��b�4��9��E< ��d��g��M�\����׬.?:�/zo��Q#�+:��'.�~�_�Żl��	�xK�g��D���=f���ܢ�:��]���#�꧖�"��@�<�Q�,+�g�����;�f�R[��l�}es&XlxVHYEB    9fc7    1fd0+���1-.���|No?��$�Q��IN���l�d��l�Q��$0�(G5�,�aE'Z��6�澩<����3�{������O�D�d��0ۣ�LP��q��0����޻����'�K���	B��.�'95��1z3��/Q�Y	�W�ꖣ2�l`%(���?������L��`�ܟ��7�!K��D��oT����~O��B�du��4�g�4�E��U���-.@v~#�_�^l\�o�|�H�4֐��^s�|^��F�^F�B�P70��;FI�Gb�G��-=j7x"��u<𶶂�s�nz�n�����P3��<����M�Qȁ�y;h�B���:;%a���p0�4����c*��b܃�G�K2[�؀,We�A��dm��pܢd����Z<t5|���Ο�{�Y.��zA<4�<Xfb�gB��Ź$*���vϻ2�'<�� ��S5^�wLg|}E�{j���z�(j��~����^=5s��R���+f���Vʸ�=�Ӕ��#�QM��5U-h�灠E�S�:ٹ,��H�:dE#|:}��۰���Da���%���5։����~�!uw�%�� �U%>t��	b�k��wf�f�I���aI�s��Ɨo����ڛ�I/�2%˶Op;��[$�B�a� ��H�d��Wܷ����ZAyΌ>ߛ�C�Ԧrřfw#�[
l�C��K^��BJ�(�m�X��[Pݢ�[��q�5�݃0~��兩U�<��q�"�	)��GB|lNOw5�$�����c��7�a=<��!v���r�p��<�o��*H�:o�]Sc=�ܫd��ŗ�p��2Z�"|(��N��sH|�L��JǫvX�ʖ5ƥd*"ǂ��9�|�{^�b���x�Hq�栞���$EO�)!?�[��v��(�3��H{����	�W�H�(^��9�G|7Ǧ��݋S�ֶ�.��.r��?��s?��1ݤ` ,������f"�ۂ<�s�>�ˏ�oxa�#���?Bc��e=�dKOH��ozo��O��Qx��%�3U֣Jz�G��[�`m�e:U2'��x�]I��REj��]]�X���o��;j�L��e���d�
9�u�<&k��rPp���u��b욲/<2a����'��y��K,�����!��i�:[Ɯ�K�= L%֨�;i(3_�t�dy����y;�#γ)ʯĩ7�-8fdeɗ�ʾ�m�<)��Ix>��ܕ�����j�_���!::[o!�\���PAr��a@T�ݼbz%`���2��j�h�JWgY��~kˌ�v��u�գ��
"�ݩ��+~lt�-J���)zv�Gq���Uh�0�m�C	<})��o*�}�P�HY�9�EnD��S��z��JU����ߥ>y� Q��������V5�_���)n��oe=�u_�1d�� �����`�'9�8?�i�;)�Z`��H�K&n�n��S:�ŷL	*7U#t��D`��N�_a�V���%��A����>��:Ja�Lʛ��r�N���C�Z���$�8�䮍�����1�@q���zB&�˖v?�7�O�p�6@���i���AP7�o4�oY��c�m,�@�ʎ�����P��U�0�*��.�w�NẬ۟���LCl�CR����ˋhO�g������t*������3��?�,X1�B�f/Α���� �$��)�;}���{=+$��L!������͠��%�=�j�$��!5��^��I��λ�Z�k�&ˑu��+��2�>;kM� C�c�*�z���N]&�~]��o%�$�����5`�ǆ��D���Rd�i�Av�#�G׆w�Fv�����	�����gL�S)*��ea���,����*(S�	l�K�Ka65�u�`e�iu�f�����%<��O6|��Ig���M�^��P��t�e�����200�*��1�X�z�`��n�1U3{q<$!�l8Ў�`���5"�61r���I��
�O�/`B�I�l�:�sҠ������%3�H����c]P�kX	wE#�6�i��	���5�P��`��O�T)8y''�&:�߼8nL�� ��Ы�h9��yth�N2�����t8��S�`w��㝮u�vG�M]reND��6�
p���CU%1R�����:}m����U"� �H4�%M������ۜq�@ya+��m<��,m_N���hf��¡�\�"�c(b���DX���X���<WwcjHN6,`��͏J�,l���bϙP�g Ɵ�?X�����f�n�# �F��%z���ט�<0��lY�F�ْyV�ͻ՟<YF��X�˥p
��7D5�Ѷ�wt�2S#ޣX�u�0�H>��M��ߘ�n�V��C��'���}������1P��xLY��;k#���ʞͿ�7r��Ι:e���s
\�p�9�~�8b�����A��5��������B��3���I:QR��gc���@��d�'o�Y��80��e��?�p8l�lmO�Ҥ@����O}�Ji���67�,U23PH;P�dԇ:�~n����0AN���̻��y��uF7=���KF�
Ya��ʃM���oV>n�vK��#�K������,���g$<I�4QFx�y���Z�tiZwe`*E�s1�/.<�rc�$�0����h7��H�:�b��B�o�"����\�ݝ�?��$�~ z�X�h�E�ڬe��gk�����7 ��3�)��r�kkX��:o�P��W�Ԋ)c���� \������<�6��g�D�K$#$A�n�|C��+�K��L8���[5��2��QC�!f��6�>$�H���l��9{ޮa�µ�]K�����LdhR�`� 6�U�]���%JT���~B���hëϹy��t0��!���j槹!����l�*ksF�+�]��5�%,�H�|�q���9��J�k���=\����IV%�pd������|�і��x��'t��%�nńrU��'��AT��;/�uż$�b2�ps�\��u��Vh���!��=�n?�+�@U����W�b�J�<I����G3�%cN��V��ܨ۝�L
�Uek$w�*�ᅊ�)�V`�7�2|��U%��+M���xo��{��+.6�n�Xa����W����GkD�F���P�c�
�� i�-}DQE[���*�~q1�`�%�)�����
�ΘBT#-�9֓w�Pm<g-x��ٰ���{H��]r =��0�Q�-\c�V��$�8,i��&�f�=q�~=���*��Mu��:f%~��
Q����ICP��B��Μ'���s�N���U����M]�*�A݌�H��D���3?�*�����O�j�D.�@�����R\&��L���eQ���M��(!j�W]eNL�TU�o�'�o�3�s9��d/��91W��_��F{�s6�Bk�񵍢-�9�˳f��a��S���hTs��<��U:�wV)��0�8i����ҏX�xu��9�/ bp�?�`����ĵu��xE���=���W;_��޶ܢΉ���P�k��r�����^�)�6��9EV>����1�/B�(Q���iS�k����*�R	���S�;�;V2Z �:|{���q��Lxt��/w���7ˬ[X�o����^e��p���8-�@'��\��#8� �zu4X�Sz���8�>�ae�:F4�����1��09�����X�H:
�������gu��gij�� �Y��r�{����O�k>���cn�o��[#�Dy�վ���@mnY{����= i��ܹ�B����/�*>��-Mb�'�H
z^
��|���d��t	C+�����t��
�v��p�@��f��eY��-�
9��g�ځjVVdy����*Z�@$"�>b��:�+dN������V����!��?�e�IK���v0������^��t���$Ur5-��9��k%�4/n�U���Lr���7U����>�2���k	����������ƍS��=jb�Ι@��J��]���h|@�M�rlT�a�O'hd<���QtI��h*�'���[��M ��[�p�Z���A�{^���%c $7쪱�T�Ep��9x$t׼V�߽�6�ҩ��/dBc�Ie�/i+Ui�ZS��p�������w��5or��R+�x���B϶�3���J�&>2 ��58��"��\,U�څ������:@�d��w��ٙ��am� �0�����E�}ѯ۬7�� ���b��n��n�ȅ��Lǡ��O��k6(+.�w��qVџH��)��`�$.� ڹ}���dݓ_�F�|�0��*�\�:�c%����Z҉+���������Fj�����8�� r��{�t�7)0��Ka�H����M�Di�5�Ɋ�u�W~��5�x�sf���������|sb(1����5���a� ���(�Y�Z't�H�1�a�K#�ٗ�5�2�j}jval�|�3T�.n��i�C͚��&g�ܓ��5�68v���R���py�`��6)*n:J���=��^CoV�}0�بnyч%���ݟT�K�!8wM� OQp�AПr#Lv[��z�R[�p
�7W�����ka�;uָHJ�=B�d��j��ѐ!�.I)�7������C��mN�&pET�P���bf~�.�wl����˕�����v��"�Ϲ���<�5,+�";�u�A��/@����L����{�D�����2�."��}̕�Gbr� �Ka��b9�F:}���]��*��9��Hf^�Ъ���ǻ����)1d�eLr����}�f�;��5��/�m5�e?\g\Z"r3�cD�����
�88	2.�% |���N�⨰%�Ϳ0^���,�n���*u)�����[p~	�7|��.�������P�{a9S*s0^�z��L)�X#6�c!2&Y(P�{n`�WMk��c�3��Pc�3�l4�jC��խ6cD�=��SG�Z6s*.�A$�E*��^�YI�eB�^Wo�X��%p�����Tu�!c��~Q�ו-
,S��}�p���A/�D姈_��!��R�wU2�KN�Q��<3Nc��6�&�O��W�6xIث�WEބ�o`���S��V=���m�׷��@B��ؕ�ef�'e1V'H���E%�#q�Au0��Ɖ�~��M:ɓ�wH��CYI�@��<Ȭ���9�Z��ݫ��jZ>׫�ց�w�!�Vܞ7X��Eh-��,ɲwi"�X�a���O��X��M��U�`-�'|k􆉸�BߵB����&L,7�Pww,�'�@�N� =sTo[=�JL||a.�YU��(������AK�m���.����کh4����7�%�p�q�"Do��6f��5��V}���sǌp�Rf�|I�K
^���o�!����xo�P������7i�%L����4jH�K�o�Es0�P�Z©uƝ�-��G����i]�8����P�m_i���v��(���k+�Y�1�����0SX>6�61X��F}KYV'WH�4�[��{r8�7���K� 4x��j YIvߏ֤v��-}�:ޒ�s�3Ep��@\n��f'�{��`P��]��´'��A}$���>��fg�r��[X���5i��'Cߥ34�2����V�:����~R�K�|��"�C�و��H��B����d�n�^ZV�PZ�h"��w�y|k_�h=�)E%��Zv�a��L����>����J��ٔ��u?Z���2�P�R�� �&;�1�R!��d��$g�M׊`S�ex{n;$,!�T5��H�}�܉��O���H��4�I ^�DH
�F�O��fy
�7�S*H��x|H�u<���d3)����캅�&�����u�5G�r�Z�7�񉞛D6��
� 9��Ha!Oi�s3/^�5��%@I��=�H������ѐLt��iQ:�5̣��$P̌W�ķ�JX�=��R�'�%6m�����2��*��v�db�]�٦8S���`,��J�TF�~tuc��
r%�X����ŏ�M���B|T�'��K�Fk��%�rR0��F�L���H�*₽��K�����_���"I�<@d�%$���ߢ�F�LBR+�zauBE���fh�����<�r��_�R�KQ��0�T�%"o����7"����A��;s��i8>�B�%ڨ_?���ȫ���!*j�u��cmd�?�aam�D^�Iɜh���r�g������:�Y��M�I��<��HRa����[��~��"�0��R,b�ty�0GP�{zyck֤�֠�5��'���tG�B��x�O���aE���������0@2�k�Y���(�8�8��H�@�-��<����W��pi�L%B5��p
�뚴hY
��a�����S���m��|V���Z8���gK��#@{�|�
�L�2���"�x
�a\V��h����������-z�?l�g���5���O4��Oz<-����.�v��1����`�{�$��e��Tz�lQ:�� �MQ��6c�q2����;,��z�XÏ�U`�x�Z�B7�ǥ�`qg���v�r�&^IMh����%����	*�Z�M�KΎ��Q�� >�*Ny*5}���� ���c"�F��p�̝�D�w>���&P��k�G�m>�3��1�j=ɇ���5o7��g;���	I��C�7�Q��k��cvD�	�T5�z��;]Z��y`�mZ�b	��p��q���t����zزP��Jܨf���*D�,B�<V(U�MH�OE���Qm<����~#����]t'}��*J�2�U;y}�:���k��p�-"��L��@ ��pA�Bk�Q<Ɩ-&E�Yb�e(MD�2����+�0����3��0�ݘl:�?}z���֠��uU\���
)��ƾE8��6Bhug�^�b9�a6�q|�E���xY���(a>2_
z�_�)9�9\�l�3d��4 !E"1�ԙ3�����3���ӧ�X�Ro�s��n^���o�X���_�9��45�,k'k744�Ŗ��ѝ��cJ��ܲ:��'L}�\�y7���	��;|O��>m���M�~w�l_������w4�T�%�b-̙�?�9S��V�>_d �°��A���t�:h�6�M�U�
�NL�R��^l�x[$�k.,CЭNwM�5)߹s　��K�I �c�_Ā�ǫ���9�:I�~� L|�C�_��Q4j�b�`���`���35��E��x5Kt�υ�z�z8ey��kA�����$rȟ���  ����ضI��%�6��B��Gε���o?��;�
@�������-L�&�"5\p�܄e���t�q	~(�l�v�1�.X����o �"�g0[Gt|6F,rJ�1P��z%�����~y��"�;���6�D?ju���|)h!%�Ŵ��vP`������U�F��'&�P���d�=�L^.����O�ќ��I�!$5'�M��7i��xUc�X��C�1Xi0}�2g&�w�)��\��alѠ�FT��_�&��)�D�q=�u�%�W�%�B�������y�l������x�a�w7�(c^���g�A�5����43�8�5]Rk�au���ͤ$�c�*��,X޹:���h#o�u�g�؉�x%����jf�W)�}�M(Ɲ�h��2�o�Ƥr�·
Jゆ@�5���U�y��Uə0���e[���y�0nO�;�[_Y:8΅L���k���$ߧ�h�	ݲ���DM�p\n/h��A�קK���[/��9��{�����d6��x�i�\�@�_hP1����\�-�s��(e�s)�qq
^��>)�5�zy��ZE&x�0iҫ�s���T%Š��
����p��{~]�~�����I-9�v�|��cV㝔c4ܑ�e������yט@�gc
��c��ڥW��~����s�qnYByٲK1̅%-������ff��ñ���tש�x�8��Pq����@�-:iq����� �5�^��֠�����k��{�