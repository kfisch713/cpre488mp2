XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~�I+��n����[n��ҧ�N��%�ìO�p�ʯT�����5YtI�yT�W
�m8�Z��4�>��ܰj��Oҡ�49k�d���_��|�_Ʒ�r��w�<T���p����!��^Y-,��-��ZG�
�U�Zn�u�����E���@OY�-�L��0u������N�����'��J��G�	I��~�3U�� ��Z. �#��U�*��b/�>��� ���G�w���a�ib	�.[�1�b��3�b+�( j��a.�6�,�uB�����h��D�(��%�t��Dr$U��Kճ�Zi�\;0B���$��(q�rUVVi� `q�,k�3G�U:�]o�"cjֹg��F�����f"�lK����C�<�$��$G����az�{���A7|gH��Z�^.e����@.\`.lw]�^��e�`pY����5?�|���x�wӆ����C��O�2����	���D;�x��t��mи@y'�/*�u)���3=�W.��Y�G6���A����N�}��vټ+�y��*S\����c�RqxY�?՞M����@>��n_���ފ�u� 	LM�[�[t���[��|���k�q{���s��N��~��g2�������g��c�ȭi����fR>�6��<1u���DNF���_n��8@`�va��ì�?7��5�u�Orj�5��7Ԋy�������.g j���Ya {�=�����Y6�q�~� Кݾi^o��W��_�v�b!�37����BDFܸ�FXlxVHYEB    5cad     f00"���������U��_��b��N�=�-j/�8G�3Ժ��_k�J_M�*nl]
v�����m�����xi���F�(D�(7��]���W׹��|,��_��+obO�G�\X?�V���8{9	꿢�G����[��YP��ö�)���[e��聨�\����軸/3��ȗeI�L�͞)AJ����Fܮ"#6n�x��U3j>�H�q�[��;��d��{]�)�ߪٸS���7^\t/k7[�G�ݽ˹p	\Kl�6�0�����!#�3��Z��8[z6��ظ����
��#��Hl���=+�?-�q�����&!"��D"��|�5�i���i���̕����芜����]`��8�Ń���<�^�OV�]y�i������y`��L|�!�[�,��OU��lYI`���HR�TC��K�U�òg�H=s���-={vjX��2�^�,tX	�
�x��4�3Z�^�03�H�[�$V�����<���I��J��c�Jj����M�"0{�4��zly�l�.��f�|J��B�R�����޸�1qA�m��Q�btrK����B�QK/ÝoR�x;
�g�y����үLm��u����M����Q�\A/et���*��kF�!^"bܬi}�F�]��+��"�Y���|�Uk(A���q?ي��Q��tN��rq���N;5�	.�O�#�o7:�S;�6�����>��n�"�!��i�F����eY��0}`2E0����0H�&��"��#Ҷ���i*:FHq�X�A� ܫ�N,&��M\þ�I���iJ?�)�gtƅ�`G����#u?Eu7���`���I�y)~	�"�@52㆓)%��,Q���ۤ�T�G�Z������۔�[��f�7?	.=�ᄖ�Yǵ`��I;9j��7�EI�,0^���|�h�`�ea�m������t��#�@�[W!�
͈@5U���´�?�8���ֻ�or�Y��t� �h�+E��0�dg��N$�H��6p���g�Bٸou�`����20v㹎�ZW�028�����P1�f��'4��L�p>p�Ծþ$Ĩ]�%�3z����-�n:"�D
e��L6��uJ����=��1�k/%��a{�bq�� �W��C�5�r���N`�ٟ
RTĭI'v�[ 1ąҢ\=�l�t.r;-t�(���n	�g7T~��]١vM��=1�����C�3���`�R5��q2��h¢�u$.v�;�J>@��W�G��o�3�q��/���b��>-�=�:G�,����Aќ@��f&E[��l���RMe�=���X1�50����Q��N�)l��%e��V�w3;��G�Jm�9�\+��hT�����K+*j7���Eqn�a��y����3we[�4��n����H
g�X}Vڕ1x^�uɅRF������4�)�B����V�a�.������k0y�;b���'b�X���ό����T�.�bf�p{� ��k�}���_���xdw��_��)�G�V}��ï�MB�1��'���@ӡ��N�I������,�'��풺�!��5�?��Cn}7]�T��z��U�X�%��W�:�zU9�qF���x0�Q��_C���%�)��[���7�1��1�Nćk���㢗�[lT���e��f?t�J���$�E���R_�k{��1)�)�%G�ס@5�^kV�z"��� ��g����o��y
���qT�%�^����;1�I@�&�2���
�j2G rB�!M��6$1�0����3v�Y3P:����8�RfB�B@(/�Ͽ���sW��������o�&��U(��@35Rҫ�����b^��/����"�뾂����ב
���&3�����SSs+�������3ݹv�4�����K�l�_���d�S��D +H��m� �'��C�� #���f�E
5KI+�t8U2b���-?;��Μ3l�ݑ�*&r�/BD��̈́��T��IA�ѷ����c�	��aܡ�h�?@"�e��:[�W5����X���QZb��si�ߦ��:c�u�4�abJS#+0�NWM߽o
�橉�/�Mpψ?#}�8�N�F[\(6�?�}�Փ{r�ª�
)�q\a��=~Db�4�=;��'c���EG�%m ��gB�'vf����}[��?����	y�;03�)b�qeׇq/�f;��=�0VP�ŏ���6)�_��5d735�~�W��A����{;��z��NԻ9�Mu����xj�?1ɔwY�!�&Y=�xk#6}�PQC>��6��PO���7���T�'ꝘܯPJ�Û�x�`׮�h~�)#��itΡy�J���1��>�&�`e�er�r�g�e�fW�@v̽�w���|�DKn�5!��l�I�=�E��P1�Cq����y����]��)6���p�@Z��N���C�>ɣJD��������x�@0��M��!ӯù_�=F�N��Ӫ8�ϾҀ�����V^��|>z�����Waș~��>�����a�y)� |߀�aN���̷��@6�[�h�����ݤ7!<R���#���)Xm�oC&I��z�eN?����M������Q���t�z��8G�1v�@�a���@o�oD�Z��&<؊?�,�&a#�@� j=�JX���>]��&o0�h���<[��^yǜ�|����;�Z���*/E'�+�B�h�R�u�+>5�k��eL)O�:u�3��F�����bW@��p,���=ukR.r��]���>M9��/�P�_�N�X����S��&�m'�a}�c4�9ģOØ[�Y�� K=��p��A��a܋ ��6�:�eo/��pQ����6"6cU���̗(��R�+>���p:�h.��
g�b$�5����$�0�8��W�͛>����zTjz�d�1�=1
2%��`s�[J���������Z['[���|�ø&�IF&�"��sY�
_^����8	նS֚[���+j�O��j0��\O͋�[.gFse,-[���&7��.*�a�����צI�E��2g"�Ta��M���`�l�mW�J� �!��vɾ)"�K3�v�l���n&JB/���ӆbl:��(d��D�dڅ����[�h�^h�s����&Mc�B�@}<�R)s��|𞎭���[�tnw�2<� N6tn+�,�'}MBK�_H/�3C�N
�[ҿ�嬓f[��5�r�A-;�5��؈�~�݃����pe�$(�b��@�ߖ����*�R�|k6������w;6k� �}��r��B���� �Y5�Ŝ~�n��х�/��K�����C~��⒕����[����W�G�0����Eh盼���
��,�*��TSS2�X�V����b)����}*[m�y�M=4�8K(�^"t�zW��w퍽(`!@�$�*�0C�ڞ_V0|�=��2��h������ |A)��5D9��͡p"�7)��u���s��W��|b�2�%*��A�őT�5�c�,�e�Sv��K�U��X�]~�*���PǇ�n7�u�����Z�B�`�m�x��$K����zB��$���k��/�B�fl�#����.�X�G*>Ӯ���\����V��7X�0h4�U'#
yE\@��*���)<��q	SJ�9'i?��YBp� A��S�٦GB���!L���{���W����k��d�K�Ob�d̠�<��FNY9��̡�ٔqdwa��c��[�{a�.�q��c�p�d������

�oD0����,���[I��KRlh��?FiAo*!N