XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���O9Y�3X��>NK�@�m�4U��������	aOA�y�D:,G+ x��L�HH�ϼDgD8S���S$9/�|��x�S��{����x�٦����g�8�q	N[��BZҌ�@"Q�}�C�n�����͢3_�%ANx���$
���;���e�$�pjt��X��`ה}h���-����#���Z�]=��A*	A�_t|oaO�~���&s�䓾��[]V�j���l��׭�<�_��٬~��w	X�/Qs��)�qp��	�"+��41v}%�p�5ik�Һ�pr/����F�1�ST��M�F)�to���$�Ǹ�.5Y�7�@pUK�e��gmB�n$e6��[�t���и��3�8\pԀԑ��`Ю2�6��*� �x�����)+[��)_]SՂ��������v,P��GCQ���%G{�g�D1���- "Sv�o3�#����^Q�'s��O9� ���.�ƣ�x_��^��P��;���=H��]褹����`���e�C�;�jC�z�d({�bN�\DF�(��dM���
ڦh�T_>�KUϞF��fH29��1A+�I<���eR@���;���A��|�!:�iW˳�����&�i*K����,�Iw�$Y�Um�◁@��T�O�U5C���8����v%��Lk��p/���'#��ɧ�&>@;G��5d���O�oBC�����	�nt�I�����>�l�-�"�΀��PXlxVHYEB    b087    2540�D�Ы��,l��N���!x�n��uK�X$�F�QmT ����GḤnL��(�[W�:�cV������@��������?��N	�B�|���Zf��h�!�k�<�#hƚ�pl��|�se�)3ЙըN�n??�Sy�p��I� G"�<�|�/v"�<ޑ����` }?�OI*ȫ�������V�3�	��5�&�b��	k�"�p��� ���1	��߀o5T�	�Yy��&�a���f����c')�~�����r+�|I
�S�I��闍��ۃ��Q+x����eY���:�R�����o3�-)����=B�c%S�X�q5��݈�W�8��8���(!����	!R$%)��9B�ّ��|$a�]t���Y"�g�UR'�3��g36lA�*�-�����,��wϔ7夘���3NC����ó���6�n��;1�S�w{
M �CW|h<��}�Kɵr��mw�."���ͫ�� *)���!'��\�NZ�����ˬ��"�υ>phm�M��Cx�S��j��0�Ͼ�NEo*�ۚ��* d�*c�����M����?KKEN�)�~�������J��k���H!�#)��t��p1&h�{v��H��[Q5i3�{b���=$� ��<s5�&�l'l��U-��묁Y�Mk������(�Q쏋�Kو�{���0>���F?�����pM�l�Rc���v7��#��<�"Z�buJLb���w5Z�T2좁���UԤ�=Wl�~�
9��c��/����㖤�g~U���ҟU&��r���I)�g]����+���~C��N����&��P��c*{��#P��7Z���C{;ta�:�	}b�2L�&U�u-�n��;�L���'�k54Μ�߂�3:q�x�� K��{�f~6��3�egG:2��B��C�{��Of�8A�Y�{eΗj���H˿R��&�P��2��~/�B%�!Р��a���_Z������?*�8�}��y���X�E\�j���y	ˬ��_�6�X$`nV�H#L����/-҇����A�{k)S�� �
]��ޗQx�,\���JB��7�-�i��L^�w������SL&�#
1>}c4!�嚈�79�ڹG���sV�����.��^G0���%����-n&la�i+
-��Y��O�ML@�ʓ�Б�j��ɇ���{��<��F^{�G`� dgqj̹�+��X���<L��˵c�� o�G-^��8�D,��ASp���KGȴ��ny�^�Y˸E�B.��ֱ��7�l�D�~{�?�^r��v�D�1 /�;f;~�'�������_�ƨ�4Rm��$�u��6��$1����5���e_��PV>��N�Ҽ�p"m �����L���N�M�g��m��7�"�i<��vg��)V�I���SՇ���u���N��"�Qv�T���r�!yK��?M��za*�,������S�P�x4�i^���Z8؂�F�
Z��U#����$۱��fc�oP�����|�(`�>_I����4�TY.B	M��ؕ�;|��[]}��y0��-w����"�	<��?=��6F�
�_�)|����Κ�{Ji��ǧ�k�<A��}�Dw�Qy4ē��s_�>ȓW���G$���2-�[�7��8�s����v��g]T�Jǫg�i7h�h�T��(���'�vLz.|��&�ϸk�Q��L�-��$j;X;�2�^��h�Wn�ۀ�-i�t��+�ֺ� �-�@H64���v����^H��&��Uj^����]x[��>�-��B�� ���F~�p�!�b��Q��r"9����hҵ�H �$Q�~�;|��0ʱ�g ahZ�2�dI��U���F�Wqt��2��J"���3&�3�j�d��Z8��,�Q��G���BLփ�1�.�]�w�82���4U����Cu֝��ʙ�k�S�����v�~K�R�x�Q�<E"��=�˦:���"���hK�"�qn��Z%id"0�T�<.��N���|�h�S����D���K��Eg�z��+�;��{�W3=�ӢNa��d�a{~K�]na��\^��Rؤ,p����];��n ��ty����,XQ�$G��ϋ�dE�%��2�-�B?��5Q�q��<��h:�tKtt��P�<�&Rf���Q��^I��H��GSLhAT[p��I�Cs��M�	C(��^{�i��<��t�N2��7A��SW�F������}�I�j��N>��C�;���O�L~d���ڶr)g9h��۫0�nԩ�X��wMW��J��nR!^�$<,C'N��j�Ax$D���U{�Š/k�9��^�&�>��9,�f����b368�<�?�B6^uϟI��)1�A��Ԁכ����C�����Q\�T�U����:�/ُ���R�÷Ȋ�܃Y7�<��Ã�0�z:�o"��9|)�
{��#��`O�~�B�p;�[��4 �>^-�G�fB+ؽ`��	P���ވrW:�������;����d>3�(�����J�7/j�ö����@���}K�h̋��s�!]F�M�8���_Z�ܟ�� i �K�,�fq�>AM��~�1 ��{k�zծ�r}	�񊁠~	�eN�5N��������Y��uqG�� ��8�ٓ�����s�D�:�>���tp)�������[��v�!���[�u|ͼxy@j��\��-�މ����$^���l֩v�5���u5όԤ��SI�Q$��Vkd��	�)�yZ@�+W_�!�N�\O}������A�,:��Dt0��D0�+`(:���T=�{Y��}#�������q/$��uլK@�3����X�������r�z����y�6�u
;��	7�3��C�*��R�E%�?����� ��۶�p
$��+��X�?�6��L���#��L��;߉Hi8��:14o��[�H%[�ߒ&�&���Y� ���9q�����8zG��]f{	�U�s[�)꽢����I�#��%촳�d�e��)uv�R���8�U>|�%��w� ����}��L��>�{�N)v�E�)G0[OF˅ ��a�i�FBt�^ަ�EqVѵ�:�}��9&����r���9:���E�U�N��E � T�p;~�4]���譴F���h&�����U�� (��Bj�FJz��r���z�d�.�z�a��X{���S�iG��|��[���h� ͐��.�I�!�t,U � ���:հn�ȿp!P��w�E��h��Ȇ݊4�U>4RϏ�PO0J;�΅ r����{��\5�;Zf�4.&����d�o"�C�{أ�f:֜7�f�e�\}�+�l�s������ę��p�y�p�^�{�@d>W�@^s� ڔdqɌ-�Z�������-�Hu���C��:�@��v\�
fN�� �~1�Km���]h1>vRv�����9I�0E����@�VF�M��
i�|ap��=��2��]�;��S�Y���C}�=���˓�2�bEz.����`]��?�x3Z�<�8zo[Ɵ5�]w`�+�֝č�4}P믯䝥��r?����^�Z�5��oyɎV�Hf�x��K�~��lZ�����vAqZT��zQ|��_EN|r��b_��Vi�!/�0�:Faƹ4{w|�7ν�� ���2�E��� =�6�1V��f��l��^�TlQ��������A���Pğ��!LƢq�zdӺ4�~�^E�*�4C�&������LLpKk��L���ɍ�6/ۨ7�6���z'&�y���`�I���ݕ��& �WȺ���p��P�ǟ0�\ �C ��q���: vQ��x.D#R�6<%���\�X�6�udrs����P�Y�a�Isz1� �m��KNf}�g�5�X{���ălЛÿ}�)I�	��3E� �H(�Y�x�:��-Ҭ���h�+�TQ �-`e]��TW��ܭ!�	u�����������!�4t�'�@��l|z�VY.טa&W�&�����@7�6ӭx���~%}cmPe#U���6��)�	�X��ea��_S�=H"�ҫc��.�4XZ��Q�x)�5��x��ւhՒw����-gZ~\6aןַ��'�(�Άa9��1:��c��OLi.��XT��)���T�\�� {��L�0�p�?��E�3b�C��^�#�Qq�pw��vpGuP�]��\��OS�u:R�<h�B
Zg�;�����V(Q�g1e{q�L{@(�&��TnU\��� �3����%l�N���kQ�#�e�όR?�B���N�ޙ���\և΂	�����NL�1)S�ʈ}�/(8�YLޤ���	;�G����A\�FA�>/���}����y����"/����!����i��[���Dȵ:�mΥ|�õ�Wr8d�P\;p��%���?.���q��5��gg�p�� �ƌd�UB��ľ3��C�V�B����2~|@C	=Ҫd���ߌ�_z��W3>��1���ag�����l;�C=��zμ�:X"��l+\�8���p�n��h0U?̬;��Ǖ����8-���)	�UeK��h>�'h(,�L����:��e7����9��ɜ�\?#%8��<�y��!�y��辺4B�I���m8��q�o�4�]'�ļ?_{�N+!U�c|�WJ ,�bў�n�]�(�[8�Y�z*͞&�q"]�F�ȳX&\�tX�$�Z�ɸ��o}x������Fg�����%|. G������/GG($-
H\;�U�i�'·~�F�#�;��J\$k;	�1�s��bZpH�'��b��n�мɝ���`�mZ���V���fQ��b4-d&OM�؃q���(a�$�low���5�m�=�-��d�u�X�s�W!h���+�5UY�����{�_� �&�E�`�	 � ǯf��c���2Dx<z_=�O���%��r�1;>/n���ԑ� +,|l� 6@��bsJcTs���W���g�	�}'K����,؅��?�zy��!����2V������ڏ�.�6S���~E�@J4
>�y$�-2��]�I�+��d�QO����� [�TN���͆T^����T��d��j�2S�O���h�*�{Y�I�6癿wA�:�A����i0�:�<!]�W��\nW�aFX���Y2k�.G��u���tA2�f����M�b��dR��
C.�|=��s�IJ�-�i;���q-�=����aԗìu���4�AH]��ْ������}�i����>��j�,6PS���Y��njr ґ���%�N�=2��cK�;~��I˚���˔c�dJ5��1��{N\H�[0�G$���#V?ʤ�ˉK�Ü�E8�+%�`/ӕ˅�M�>nY4x��q��dN{��S
�)��\�V!W�0�Җ�<�>E�Z`8{�A"�ڦ��2���Z%.��B�K�K,W�k*{�>�H}�mw�� +��ATR�RL����o"�^���J;�01u��m.~n��*�j��v�x\�CŜ����nL�e�OG�$�g<5��=��K�ƌpxW�d��t�������9����Wݣt=IC�Ԃ�cb {���IX�%��ա�#v��2q��k?5���!Ԁ>z�������r~��a�qP!����CD1a�n9����E�SJb����m�ꁪ��u��u,*bl#U�����P4�e����dG�;n�����3y|娚�7�[�F��Έ����c����ɕ�(b����s	������?���R*�u��V��
�,�,��͏��Hn��P���
�U��s܊���	axێm��P@�$i�M�y���br�`BJ��`�O�|��c��#�ɟ�c�p��I�P����$\��uF��mPkL�(�)�*�ԋZ����#ff�MB)ca�	w�qIM�Y)0\���CZ��`N��8TI�]�d����@��ւR�������T��e|������Y��?��x~}�.���',a�/xt���c@qK�2�iW0��F��)��O�b����ܟ��V�c��!��$̥��3�y�f����47N ��.����,U��zX�6�T]J8��4�%o���cG���im��zv��t�X�)�&v&�7_��r>�s��X����n�̤Eվ����δk!)�g'b%5�tu�U�x�;�����8��R�,��h*����lo��ۍ/��J��O��5�qю(*cK�-����.���+�)&��{���L��@�"Jdc�J�U���r��}H�)_�2G�*�8�f#��]�E��e%����J�vg*�a`��.�'�9�kg�V��Ņtt��MX��f��4*�uR���c<Ȃe>'�@�ƺ}�2���i�n�B�J��f�7�-��M���\�*�G:˼��h`���=mA�Ӓz�t�̀H1��b�B��f�������~;<&Qnmߠ:BE�w��{�K��B�0�h5|h��Ŝ�y��O<�dm�D;���K�!����O�B�*v}ni��؝jZy�L+~c�Q0lY̾�4��mΖя���#�o�����0}m߳]�[��v(Z$G��|�ɓ��Ɩ��s�3�0��Em���0�dZ�+�zvw�B�`9��0:�v*MKX����MH1�.yH4!�Ԩ97��"%�D�@�+~���cFPe��"���(�����"�=?��=	-�쑥D�="�xk�7�-�����-��ef�/��zf;��tˆ͆��Ť֫q|��f�˽o��3��-�(Кx_�op}Ud���<�9��D�d��5}��=!�R��=��@x���e�!�̭Kl�C\Li
:�Dy/�I�� ��;�d7��Ƴq7�) ��(K^Gr��oƑ�%B7�T�s�@�{��>��Q+��������c)���GD�$�/u�yF�-ÕOc��n�F��j��>ε�Ȟ�W�@~���+o}}0N��_�G����Y�.�p�Ԡ�*$��g��?÷�=� i �@z�UE6��/$=�o�~�&�o7w��w�sg=!��Ϧլ���У�%7��c�	��3����j���㵭n?�M�vZ�2a\iAeL�%�W%E%?�^�������O1GN����ɮ�'��_D��[�+�ϳ@��7T� ��)v*V:'���b:��%��c�^T��S��Cńfm�+j8�����y��
�a��Yq�X�֙)��C�4��"d��.K������;�j��/��N�8ۛ��+Fݰ�����b���O�^ͣ����Ґdi��3$�.����G��f�R��H�5i\�: �J�w!���p|��o������تR�b���r��C����aKn��P �oʋ�K�` BY��a�7�D���
���J9e�mwV�������+[�cC��8u>L��ω�1Ɯ�I}���By��Ţ�˝'P2��8���뎙7c�֊�Ό�'������Ow;N��u��x!�����j�U�۵~a�8�X�k�~�=B�N�H$�<�S�L��6��R�$M9��"��"=,G?��j1��@	��4�	�-o�v�_���0���	���9��I�:�h*����ڱ�XV�w����|�ښL�0]7��^�ʀ�L��� �;�'�#�����@e���������rL�h� �K����C���������U�Y��{� u���o&�i���e��Z3k��5 	+�!R���8Õ*��8���F�M� ��Of�����D��e\t��,������� g,����M�Qp��c�a�7!��̆��a"{h�� p�ZѨṼ�2�U�%�&x��e��8��$�|���	(���4�Dc9����73�����(X8�Z8��?G@P�A���G��,��]
C���_&�Ź�5��V>�:���k �^�y'@���^U����=5��P�'��RΠ~R`�(���u�;��Q��9I�Rܔ�������&39�a0� `4�}09���W��y�2t�4b!���6-�ܫ�e/.�-�@>[�Y��*����2��d����3��\�Y�p��ԓk�}��H�nVy��i4��ᩞT/.2q�F{ �(�p@��}����P�C����4�A�Ub�N>�(�OK�5�<�y5J�F����)�b-.�@�i�\�Ƣ«%�*�9�x)�Im\.)��"��փi%RO�藆%ׂı�܁��NW��?��q$G`�o���ZZ˄�NV@��/��|7��~{�I�L)�́5RI9���0l	�����@p#�#�gW'����/n6��Ya0å̈ K��)ނ�
����>�b�I8�G���4%t>R��4����
-��Pq��M|sf]Y���HV���`�c�k �F�TPƫ92��ب0��n��(3l���a��Zg���q(���b�H�<�)����^�2
��M�����$��K>cu�h����������� ��� �XC�+]��st)5�j�Ҙ�>�G�Z��f�G���c$m�Q�̜�Z����d *���kؕ7z�x �|��rJ�	�fQ�P��s�x�[�љ�#��`�d����N�9!��*���sAb���71�3��������A�E�F15�(.� ��~�D+��s��c��&���M�8~f��zg������_�5�v�r����:�m�?���E~U��I���c���[�poLv8�&y�+�dP���",24.*=���w�/	��a:���^�Wf�����r�4V�6�wO�
z�ywea,��� R$|y�݋����^x���:YaЇ>��U�+c��3�Kc�3%�A}\��ݜn����^\�)���jٙF�;"Q��=��<"�F�y6#�ˬ=P�f����<R|"�b�o r����bE��|���P����3���m�.�Q��M�J��@ٻ\�5���/ߜ�D��8̕��t��"����Sܛ��-.h �t�O<<�G�t�b�P����$��#[�p�9����#�>-Y��؃%��zl������"wSo���'7�����`�\5S�3 q[�.��-׉�_OV,�)��n1���-���)��S'���?�4k�c�*����hɵl>�̬����,]�.�0"�4삖/��,�=����_��|O�ʅ��
%T�i�Xu��x�Z�+��d���&T�^�T�J�I�H��du|Ŭ]N�}����εsF�6�%K��U�;�,�U"XX&��V��o�V�+��� �!��Yȸ�	�f>�C5k����;�h�6�)�R�R����d�$@����ۣC�X��C�Ux*�KQ��a�r.����3f\��sek	�W��2+!�&dV��*���e~1��0r�D'Vk��cM�L �>;��>��G���I'�\���={��