XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���U�P��л���r]8�1;�-z���#i�R�>Vmr��^uz�O��g9����I<�bP��evl�O���kR�a���f_\�(^���� /��P|[�;4��)��JֿI[�٬ѓF�<��N��|�LI����-�,A��0�����*�������܇��1��M��=ؤ��7�[����(gO����|ֻ���fp�I&ih�3���.Z�w���f�r��̋�~�4T�Z�S{H|.W��w�[������+���?�hQ#\}�R�j�f5m�����~��ت���v�X�&��u�Vč�~�A�F��*�,�wy�χ������}?�CC�1�nE�D��C2j��_@�)�B!X�a
SK���҇Es�����c�_�j4y�l����Ί��?kI��2òC������:y
��-e�pj�w,�,
B�ʟ���V]/��.��n��W�����e�2�ۇ�L!9[��<s��xKz�R�a!��E���-���i�)��Ӱ��ǹ"�m����1�*�J�����[����1��Sv$Z��;_L�ת��A��ie<��Y�����Z��'�;o���?T��-혀�R6gj��O��]Fr�K���F���] ��Ɖ֐��w Z��Iza�����m[o/Db���ka�R�)�\2�8�(����X)$gV��z>j�����EQo��X�S�xx�hz���������>'��#~�7�y�
�A3�^��<����) �"�����$0u`��0XlxVHYEB    fa00    2a40F���]���G?��6o��eȧ���=6���ֶWB��@K��z~�G��'�`̺HRΆ!�J�c����|�TO���u�;V���A�r�{�_�'�1��+	�	���ML[^E7�r'�_ͦ���(F��L��쫎����fV�N�C(,P�7��b�.�
�����K^��n�w���J��4�J����ˮI�w�lGj�
h���U������̦ߚ��ӵJ��)F���:f��D)b�/[�o�|j)����%�uO���_���WnTV�CH3S��^��	f�����2̵j������_���C�x=b����u���eoacK>q��wZ��(t#���Ô���������`�E�$�PBwO�ܿ:V��L �Hjc��G���e���,�6�����k��1��O�:�g�T@�v:$�}&��rաڐjP����j̚����P�?ɥO@�|��v� G��E���2�5@���R6�S&��S��m�l\.A�d×M�I295ƽq�d��8���V<�D��.�9�q��$��u���ං�:�����w�R?H�6[R.����nn)�m��P����;z��~���''&��t}hgyO��L� ufhc����\�qo���P�Wg�ɜ�-HC\
���b��/�� ba����2��<�pZ$��0��r��j��Ne��K͔�%j���H���L��u��9��Ǉ�<�
���2��|%�4�]���?����sV�GM0�{��(_da+2�o�7pz�m��ښ2N��ed���
��V����D8qWt��"�s;��ڷ�)��]���K9¶5��5'��Dx���Jo砯���;#NC���؋Ri�	J���aM�����*	�A� �.��H�3s�Y��b`p�~�7��,e��g�V�0����M�G ��lW�1	���n���a�-�^���I�~�&I���t ������Nq��vST�ĉ�
��oq��BKs>����(��8�epziY�%��p4/�X86Ћr�u�����Aw������ {̘�
-99k��x����j��m���;M���1]?�pP�`d�0� R�Q�F�
V�4��eB�|�����,�Q3.ʇ�>�����w�x�]�m�U5r�Bps�Pкl��+�4��"�c(��ڍA�j�T\^Ö{s�hA3sp1��lU?��=Ґ��z�	$��e�8�eI�-�~9���R�D��Ē�{�m�#�8��2;op}0�3��<w?椔����y���3�.54���G<p��]�Pk�F����Ɵ>��" N=YV�
�T�O7�f�-�O~���I{�l[0�4"��3ŧ����O�L��(i
N��l�����/M��c�ow�ʭf`��V�y%8궝��1*������g������������%��+�%f�"��_��h��!�&1�i��m �%��p*�^%��UK�,ܱ`�����9�)�[�2����	���
��G�U���f��莥���y� ழ�}�l����C����K�;�۔?|�Ǝ, \Y���������F�����q��A0̿x�m�f��5������Gu��d|U���6� ��5w��T72�k�|?�"~���G@vU	��C����bɈ��q��eD��˭��|;��~��4�Zr%���y/����k�f�x�~{�/dR7��]�i�ð���J�ҩ�z/�q;�z͐�-�M�k^β��͆y�O�.e���BO��	��5��x:�֯�����FP+�X�Pw�x��z4غ$��Tqͤ��Kp'��FL��V�{����D�r�g��C�1�b��g�����#;���,.��ЛuG*uFv�T��[C���9U�g��x:j���xW���<�oUFȼ��ʧ��Hk��z���
To�*^���,�H�Ȑ��]YL����(��<|�_/$�/���c�eG3����Xv�TmpM��VN�'E�����p9����H�'�&En����s%�M�׆J�4��܄9��v"Ď�ՙRlg7B����1i~����������'dF��S�8��e��H��:-���"�'bH'��@��!�U&S��=�9��q�� Z�`����2���5�q�yT�a ��}v�1�+8)�|�f G�L�K���;��~bfZ<�ze��[JK�AA�9����fF`�X�Ĩ� �Zϳu/�Z���9�O�i��-TG���*�S�u
�$�j�bu��+-�R��0%g8�y�w0�*�\�Z�A�)��3��B�K���8;�� �;�kg?~���h�3�S��dY�_/uo�yj}Ƥ�A�C�j��UC
*-��7Z�-��"dI1���EA��t�%M�\8����޼��;[���b&��^_�p���a�����2�0& ���UR����Meγ�����u=s��b���҆��VNU5��wEQ�;�`ӑ,;���/2�-��0n"-[�Z��m!����#�eW����dBg�|���ݛ�i�� ^i�$"S�0=�'�R ���,F�t�P�[/q�ZY��$�:u�U�W���>��w[�,��U}�*�����ޤs�h�t���Z�h����[��Ģ��pM&8@��Ԍ��ĀQk�&�$�k�X��i�R�d���?B�o�W�Q4F�jN��{:b��y��K%L�QrP�w��Jg\W�-^�W��)��޿��/��cUR�*�n�F�B��󗢘�k ���:E<���[��^�Y�'�ן}�Ѥc��j� �]�w�=�f��U��XW�7�Z3��7t��mA�l��܎4#_�Jx��4�1����~R�0%��B�:W:ʆ7�'�n�Yn�X�v#�����EC8��-��Q	#ؚ^��D�t ���F�%��(*�]a_Hk*i������ߎr+:�篑�!p��/.v$BiK��1E���mA,%�V+�������������0���`s��=�I"�?�$���Ñ�D��lGGZ�$G�Sdg{�0Ă�tߐ�vsV���l�g����1�`>8m��Ԋ���	b���6�ZKW[��u���ۖ[��l&X[��&D�+�+��yA��bsź�5⟨��Ք���殡�>�v�R�E�s����N��I<م(�"A��g"���wh�X�x�f���LA�`M.�s��$�Q������\k��}��Æ�A(:깡�'nm�0E�_	����*+F�a*�%-��R �
�^�L�Jov��|Uy�������dj
�!�9 �"al�F����VOf���U��,�}Ť�I��HI_�*I ��.�?L�jp�;�H>�9?���æ��=�}T��nV�K�>W�^!��!�!ڝ*X�?)�=�x���Ǝ�z�9���r)�3B?��ww9y�R� b:���8�F2?��cMH��ZW$\nFoW؏5EE�#������Rh��N�_�_�"C���$�fuT�S9�2��6hs�/��Q�E��}ߘ�s4Qq-��rHy�aw��hXt��^�_�88�������pP�#v����,&=����ȷ��K��hbL�)4%���<�����+�Z;�*�){Dޓ���;��>ϝ��HH��m, �?�
]	�J��2��z*�u���Yvd-l�[A%��j�F���	͠��{���iP�R�6d,c���gB O�ѝu��+a���^�ݗ84�B`p�����J�>�e ]��ڻ
D^��h��њ�II��HGu^��������v��xs�\�чYW��"َ����6⠗cb�="�=�7���l��: �%�X!��񉦒͒W��zW��p�c�"�Y���,���K)�d3VfOh#Hߡ}��5�K18\ӥ�V�B{@GU�*Q�q�F�#G90�@�]){��)��Mf1�Shb�����mBpq���$��%$�~�=U1�\aW����C,�s�;�}l�X�.&�ъ8������VK��|�-�i�O��9 �()IK�x���(&�x7�%�s�JQ����䤏TؠT��rW��R T�~�B'p��� ]I��KMw�Rp��as�xDPo�v���)��t;4�u�Dy�@����<���FG���y+XJl ��Pu�fA個�]J��L���^�=�����R~3�A�	"�#�ʐ�|�?����@��p��4����{�eF�o���F���Q&��.��Y�	�5u��Zf�qM�2��-{u����Gg��k:��(�vAb�_�u�=���U�}��=�y�^���*OS�r4�L��Xjp>�����.�/�1;>��=;dA���"Rk5�a�3����i�9�������B}����o(z>���'G
9�&9�%1�P�]�^�D0����[�en�;��� p#ynug�<��l�-��c|nlП�����TvtȓF5e/"��E�U�
�.R�p��+=�dB���lm_�s#��*��̱BP#�Z����3�}��2KR��oW�ٜ&h|����)���8�ل<��I]��y�?ڐ�k�Y�!�C{9<�o���>�l�*�ْ���F�����B�Z�qg��y�xJ����C}*5r6�ű�w��l�@s�M�qP�;Z�ʪ������$>�}�|:�M�e�<%��\�Ywe4�ǆ��`�߳	�"ߖ㹤v��%���	8u�]WDJ���f봅�:��w��$�^�_z���C�ؼ�N�F
J��s�`��CԴRg��	ܼP���e;��~!i��fT�Kt�����.����Ej�Ɠl_�z�*vk�*>��m��Z�K���� Cj��řm��ֻw� �u+o7lY��(�NNF�j4�HZ\�$�O��@�P���|뙛l���D��x��:㈥u�>�y��Rn��<��Y0x���.c�Cu+�l�M�n$��g�=0!AC��ݯ�kȸ�K�Y���=�ļ�넦�i(�6���w(��7�(�Q��e�?���n���RMI�*v���YOGU@uQ�5>�N�4~>9m���(�
Y*�\�,�)m�*�h0aA3Bi���A7Y�5b�<I~�&-1�� ௖h7��~ �C��S���!�HՍَ��j���묇���d�WGƟOs�;q�MV���z�����>�j��8I{�s|����$�Y�ʑ��`4`] �o���o��Wt�t�3.n���~9NȋI��U�j�2Ob
9�$��x�=I����}n�Z��x����wp��3�t���� �*8�*�',��Y�Q�9"څ6TP@<'w�/^�T�D<T!�}YT�F/4>��}�i���ևD���\�D�k�xa��W9�%f�H,Z�\�ϰhV!I��s��q��kuķ�
�{��U����7O��,}�8�3����2&4�<�p��a���<Y��˪��|}vs�AY�����|��fN��u�^��-J��ݱF�*�R{H����)�# �r�o�w�bx�B��yk7אs]���OΘٔ��<���x�$��3CC�a���ƭ岾��D�������L�2O��j� 8L����ꚬ~a=���8~���9��h��Ǖj��,7'p�\"��%/���/����#ԡh���3�fU�Z��G�	܎�҇���@�H��sD2
�����F@Sk�v�9�������f���u��B���"��2����3w?.�:r4�ۼ�4rt��,ƈ��K���R_�Ï["q��K��V��ϱF%sE8���!C����ץ�O��^�f+�<-��\�BB��Vv[:zխ�?LT�N0�sq3��5lNSE5h���������m�s��$Yu'PׂBҠ�K.	������%���~f�J��6�x��-&�̠(p�a�_l�gk�R�{�$:�?�]q�Z�3�rH�,��aI����Z��<��|G5�b��J����>��4�����?�:W��H\Ɉ�.�I��z�6�-4�,�)�̵A|S��[�h�a���&���0����4�k�TF�T7z�_(�d�7/��w�!�F���ڱ6�Lcv8�6��	\@f�l�7e4VH��rVg��rz,V�x�#C�! Di���6}�y{�\?�4�Z��?"�P�'��L}d2��/s�@�l�/lӔ��G`�B\/��3Z�>�y����S3>�INL"�9�p�[Yu��|r����I@��hf�/`�G^\!"wOlF���o��u \"i�4<,�����9���o�?N�X�k��)�JI�������5]6�=����bg,�����S
�ݍ��}��\�A�w�i��*;ƫ����^����aӷ���)j�C����&���2�ܺ]��7|�O$�4F��#�`��+#�1!���Q��1M.���Nz������n��nH
yd����2��5��OGI���|E$�Re��� a�DVK~���2���{�<��<	٥�3J�T�fS��ew� /�'(�V�+��8|�p5��lS���T�>ɜ�a�i����u�� 6پt�l��#�F�ħ��Hm,W�/d�:�זFQ0�v����>�,������8<��|�C�����oAҙ���-z��P������أ�`)P|�s��z�>���N����nж^E�e���}1�W���_�� 0Y�sB=T1~b�΂A�o����ۜ�`�2RA�Lz����ʥ~�IU�e��Nt�jd�����^������e��?�H�ޚ{$^Es�s"a�	�I��Kh�c���`Ql".����v�=.���\ѐ9@�hS�PZ{%f����hPc��<�����-����g�5.\�P�M�\U���%��A]R~��*5��E(θaǬ�6~��������XAP���ef����9Hs>Oˌ����ttv��BB�\P|@_޾�����l���;��E�r
�廥bHԉ$#�G�ro�jO�_C�z�����*U�]�1v�xӱ��'�+w�&��0��A�J���)���ZsİH�Ry{;0V"Lf�ʌ��.rw�o��3��'�����2P�o����p#���C����!���u[�����UUF.>Y�U`-�ʄ̔4"�t��:��؊�?ø}�s��-0�S�Pn�����
k�C��B'¸��ڰ��Tp~�P�ĩ���0��z��g$�;:�W|eH^�ɮe����>�-~���<���>b,(���:w���ī���5RE*z���/�p��ڐ�3��6�m�TZ��B��h�o�oQ�Oi�����K�<���_,�������A���ꏴ�vy{$�;b�wO�ULT[Ŭi�� 1�����(��Ǜ��b{ʏ��ԏ�!����r��߈'�"�!8!"(:g�����B��X�C���c��w�I5���w�w��Շ���Nrۃp�b����n�k�x$��G�}���Hs���8|�W$��^��,.�5d���</�1�E�,�u�TJ~9�&gU2������e�=�����>M�^�*5��j)���8rz@����j�Hl Q��Kt>�VsNV�@�0P�"o͇UP/�^�7�Աf��F��'�$�|f=�"�i� �������]����zƃ�B���W9�n��Χ���<��Z���F��di�-��8ApP�[��zN����cx�*�������E%�5�ѐ�݁n)�
[����bL')���
'cq��7��[�����&�SD#>V�y��VRq�݊�L����g����K�J��o�ɒj%%+��<�9^ؼ��u�g����%��f[?��յ$c��@3=�EW�9�'�w���H��*����&��B��~j1zΖ$�����R�ۇՅ���E��`Z_�W���e鮦7tV���ļ���Ib�_�i�)���abQ�{����[��O��\5%��]�._w�^S�`s]|�A; (*y�ණ�>T�,<ܲ�լ����5G@H�|��^�������m����e B,)�����v�F%:����_WҶ(��fZK�y��JN��{�)�7p�|���l�V��r3�Pe\�y��ƴ�����c[]aVA�d��dPrm�kR�~}���\).����M]���)�=�V,D�*��Drs?i�8�EOS�oN����,�G
,���-$?�h������!���0E>6��+��	Bӟ�� �A��Է"�&����g��S�UdH^�hXR�����?E���U�d�^ͯ����φ)(4��Ǌ.�ۙE����� l�|R�N�rp��뼳�1��I�hu}�/y	5	RC;����_#w��X^�;Q6!��/J�5�����j_��>��݇m�7�/���$�@W�,~(ss�:2i]��W��a�z�T"e�q$��e$�3������L���V~���\�(���2
.�MI���ZB��������u^ݑF�,�u��qc�
��-����E~�`e܁]H[�
�B?���xq0�.~+El��9�U0�hZ���QL��3�n#x���5t#�F��t���X���&��?�I��Z��U>�.��e礐
88�'¦��5 �
SP�P�i�=g�4��$���)	�1T��������<VJ�k5��o(��rHk��{����@������M�H��ej��ѭ�@����ǁ��O�	�*&�J��,{�U@ɗL�>O����ƹ�{���$�ŁW�p�����C]�,��n�3� �N�C�U��SWU2>r����ض�BB�m�dHkH����mӚ�[����1�Y��Nh��	��{}��P_��)_p�Xs�u+X֏g� ܊Y�6+��C��������*�%r����-�t�����{��d��e��/�D��7-��dk�v���]#%��O�"�/v�d��+�=@l	ar�0�'�Iݙɒ��>�FMh�0Ȟ�nšӃw�zn_�
6`*�BQ�n+�Q�w�A�G��Jh:�~������JQ���I\xO����u!$����V���S!i��'�l�cyv���1��h�y>�+�z�c!�0���e�[V�6(�����=oHot��d�o��k�ש��������=f|�L��f�d�,��L؍�q����?��+�'���Pw	�Wɕ�!۫���w�d-��������z��>�`FQ�:K��w���5�x�� ���=u���,��dh�r���a��dk4�oh4d �|�ۋY�i�5'�F�b�薣
�+z�_x&&�	��M�W �'�B,i���E-��ψ���܀GWA����򽦹۱x���V)$82�w���˞N/`A9��ϾF��ݓ�w�����ӿã{u^0�̀�pe D��9�\G����tC�2���������e��Z�(0�3�[;p�A�ݖ���vo�7��w,	��tõ�dVh���\��=�a6���\������qq�?Er
�ur�e�y�_���%���r��!��jc-�$�������S�'ْɷРwb��vSb�^1J�^V�@��}Jl�j�:�%���;����j�����hXF@������q��_B'E�B0R��g��a��L�kx(�BQ�	*�G�����7�.A��a��?C�'��j���5\����B��]]
&���*��^�Z����3���gė�p/]+8��?F�0�bt��0M��)�Ϣ��{@��5&;%��B��.�8\�m�xHN�eIZ�f]%xxc��N<����nj��7Nf'�:tR9��E�'�>�"�,dFD~ʩ����2Ol��W��zѐ��ڦd��D��>ow�,W m���ς��ʽ�+�i,V��-+>���MR�)E�U�]1����(Mu���\}�bB*��8�}��>$0��Y>+�����T3pB1>f�A�]����R�:܃6OQ���YN�l�z�O؂5���)�?��dM)E���pc�w�W�N�� ڽ'QyC�x ����f�����t�<��	Ig�!�p��QD,.�|k�f��Hd��?��ۿn,�.�9�/�NY������j�{SQ<��-΀ӎ����(���Qs��/J[�EBHyBL����!����j�0'N#�=�6�D��"B_�KnL�a���n�b���:;�K�Q�{R~�KS��O�:~߿�u�C�7m�7�u�aAp�^���Ï�w���s�;D�	�xo$\�H��"��?)�^$_v�uO�ۙ��AT�Ei���U�oM�=��O�H&c0�x
h�F.�Q�@W��/�*bT03����ihI���o��f���mT3��7�@!�0�zm�����Qc���>wQ�� �KT<\y���mj���6��#��\""f�|xXw�N������S�)E��Xx�>R/{��R�!n�>�-�3�t��{8;h�6S�ߠ�R�����9�F	j9�2�N���8�"C>��yԷ�tG]�S��r��#�w�ۥ�>��_�P���2 �2��*����g���?�%!�Z}D��,Ϋ�pzq�����ҫ�+ic��M���B��+	��Y�q�s��Wc ~�J<�Oˍf�����"�<0G�1�,2�Sa�Ea��9"��������KOF�'9�F�]eO���+��f%�R=�H!m��Ff%=�JZ�XlxVHYEB    fa00     8e0Ќ�HH:ep�3��Vh0ɩ1j%M��	`-;x�lm{�i�/�2��7��qN{Y��b��JFIy{V	}��l۞%]������x/��LŨ��Z$�J'�*�֪����mQ�Ιq�ᨔ:{n��A����o�^ѐM���I"�Pd�-���#FT�A�)*�>�s�o.ZYDSV2�şsچ7��0?���W��a�k9�2a�M��$ID���$v�e��nI��jm߷��x6}�"��N����e��Q���r)���D�)�����tc懀������{Z��=��qEuj���U��Q��3�^�k?�,�t/e�T`�W b�CFg(��N`Ό��O/2� 	����o9)�!"�q� r��+*_{8�~5�US#�Nx%�쓔���,��n�����ϵb ���z�d�0t�f����
O���,,�����c���M0�[k\����<w��ݠUķ��D�A��@�'��PK�a�Ɲ�
�|�i��I�]��K������q��M�I����4��:g�
�	�DɅ�N���a�`sA*2���y��l�*�M�������!`B�|�����+��AR`��L��ˋ���%5��Jz#��/�[b��{G�I1���C��<��J ��S�� ΢�9ٵ�;2�N�f7:��8x��y�`Օ�FF�)vK�4d��I��]��n����1{t"��z�oϑI�j�}X���Ƥ?$UJ�ȒF�3�	��/���&�	P�F�F�8�o�l�>�a�.�6�L2�í�ϋ���fIC5j�+��i08ݸ+�=u�҂O�_����DN֤nC��Kj��F�Uj���y�81a�`'=��!����x&Îʛ�.`�Now>�SE�ߖ��F��K�vȋۼ���T���u,��a�ߔL��|��=�E&Fr]�~|�J����M�[�!;��!���29K��"A`�����b�cD�"�U�u��`�G�(����Q$~�2.�����R����B������ �l�4wa��}Z}�-A|��q�y(�Q8`�۾C���4�p-0+����֚���>��B����St_�G���i]�Z��/�.�P{j���5�@<]���=�v*�7,8�Ȟv��Ԋƽ���(e!dya�/+1{(-�e�Ϫ�]��x��"=��M��D��A�A�6n�%c�&1L24]�píhW`GT��!�#�@�p�	�B�`H Hc�%��A������F���:����#�Y���+l�&o��g�f8�g��*�,�V΂S`�I���ϙnaTLY�cq�Į�ȋ��4�͖eLS�u��-vh��^�h�2l�\H�+%N7Sy��4a6��^r�W��[�$���ku��_ 2�+���Pؿ�vᶥ���e�CC=�zx�|�`�}_7]I�S���w��4��e�����A�B�݌�rcC�aF?AΘ'�& �;n����.-�M��b�DR�r��ht���A���}�n�Ж��?m]�u��'�[8^��G�[���Q����19�͇�P� �+佞�`G����2��� -�Y�K,]��B��L�Xz��'�7[�?�>.�~~w��u#��W��/T���ߘ��8�m���v����(6al���d�h3ԏHD�pqT�g�^��͟/j|�P>�N�;=�c�$�'8>�<��5[�\�0!�\OD��%[�n�@>n�!�	��q��M��v��1�!��P��٦9�yW���Я�޽^��j�����*��B3QqMG�q	�� �)j"*�d0?���ȥ��u�3>lM�e�^�lit{Ru�
b~��B�f�i`S�X�9ò_DIF� ������j��B��_K�fn�Dk�3�ã�y�z�6�,��e��E���G�D���dQ�i��u~������G�&1Jk�޵C�K��}~	�o���(f��K*.ݮ�~�?h��A���a���׈!�o.}����
�iN<��Sa"A� t/����ɫ���y��<^�ey�0$"�¿>ȇ$
n� kj֒uecw>Ep_j��t/�5eg~}Kt��5���"�V��#�D�O����c�g�+!�E�*V3���fQ L]VĦ7��|K�<�-m��_�w�잛�W���7��p�5�l@��n��4,8x��+I����!����ڑ��0G��86t.aoҌ5)F�T*��E|Y�k�=6-�2����t�>|j��
�ܖ?m���EoY	��-����XX��JH��MJR��#c�XlxVHYEB    fa00    1110d�%�%(��qQK��F�{3�����������?RX����,�B�Έ��w���]򍐐�r�$6�*Ua��&�5A��Q���n�<���"��}��z$G����Mt�iE-D��c�܈)���Al>q��5C9�e?�������qc]N|u��6@�s׿�^�%�u��W�i�&n\��_��|�H��q��yJ�\Gd���+n�\P�Glߊ�?��(��< R�J�|�H�}B��e?��+���$a�U�^�ܰ�z�@��ޠ�0� m�^C�SN�M3֬5�b�q �e3�.w#�}�0��e�6��NqbIR��� �5��r�N�Qz�_4b�G�̭�Ca��A|� ¿l�g1Ƀ~�D�`������R��PU��Gez0�W0n�Nl���<�un;_ ���Q�C������BM����c���`\��7�U�*��4�i�t��k4kqBg��<�C\�U��1Z�g����Q��~��M(����ns��$ۆĶ_�\"�3I(6{�F���_��������0��N�?�7�d�.E�x`��:f)�5���Tka���P(�}�O;��]
����c��h�X�gW��5=Z���tC�����p�-�	ـDC�	^QOiL�i��!3�*;HѮ�N2wV�f6ݢ�J�N4-3�6�b���ӭ,���9�tME���k1�e#�^}�?@��rp>�B��u��p�~�B��ݏ��{�ů;�3s2�të�KuEc��Z.LfI�V{K�aa�w�y���[���`:�IX�MV��f�����{�K��o��(%nXl����Y�#�8�t����R�0������/��������h;=j���ο��&�����IK��o�o��Ƞ�8��O� n9z/�ev�u>�>+�,O�?&0[�<K$q[4�|��d��~�oZ����!O
�ʅ�����K���0�{��?�Lb�.��?���I��A@r��d'I����n�~0��z>?_(3��3�^6�g*��R]���A��u�p�k��4������2���f>�umȪ����U���!�4/�6acG7.=�X�.|�i�Xp��y\x:j
�Մ^j?p=�'fcHX\����H@�b�jd�̇Å�ߜ��@���-�ۋ �
KC�L������XM�V�[���RL:��*)<ns"�G= ����Yk�+V�&�H�	`JKK��J�����,>��f�I~.�%���c���|��(�^��D,��L���"��<���0�Aqm;%���>z-?V����Ѡ�Bw�8Ϡ��6��$?�<h�l�֡f��hEl";o�+�*Ų~��ǯ;SC�c�+��"��/?"k������mG�0�;Sc:����e~�@(����>�]�봟��l��8�9��&�28���`�?��0�J6�;��7|�D*?�Q�v�lI��K9��C%/&zz+2�̗t��.���xґa�u��.]`c@}.�R!� �2g
O�<���!mQ��`Q�ź1a�M, � ]���e�]3¼�ae-	AM	�W��Ꮆ���ܽ�$D5xV�(���u�o�~���e)ڣo��� ��E;ŵ�\RY$|�`���k�Ǚ*�(KJ���	0=O?�Θ4�>���	��`���@�l%�?��{:9���CG\<���5��+����<��
�Kt�p����(�y�?����N�oLT���vQ�	��C:�S��|�Bpn��׍}��P2�a=}G4`K�w{g����S��Ԣ8����#(��`�
i���,6�5��-�5��S	��@�զ�
�&����IEE;��]�vkUV<�<fQ���`�Uw��-�~��B=ʦl�$ȥ�:�����t]A�y���hS�|!��x�W!+ ��Z���J"�y"f���$h$2UX����~����_VP��& �ɣ��w�t|�W��,̶6M���!��ߖ�i��d$��������L+��A�	@d��>h��F3�FUDAS��P��&��e��%mo(*�_	|�`QZ����z m�!�2\)������}f�閁~�Mzⅵ�Tzx� ��B�=�Ĝ��P�BJ����W�ݮk�2�¸k�M'�$]緑�l��Cc[�h���~���Hx��kCWq���[u�A�| Z��lZq���X����}��ݪ]�[eʡ|F�[��ȝ��;O����]��RԄ�\�ʚ�XVK�#����&�ZD&�R3�B��no1���?�|�/ބ���O���K��H1 tU���a�,�۞�Ա�2�mb��:�!G�&�y��!7B�xP.�%Y��="�K��yWm��7n��9Fb�c�A1��BL����%Oس�4����`	���8��)J�e:�px#k�p����Bb�!�o%�����f$h�p)`b�p�n��c����e1����ge�5�kP5<��^�����9+"���:!��1��W�)�l�*("�[��,�~��(�Y�+�0:�Qt{�E�Ї"���`%��]2i !�'F"��F��|�)��e���}%a���)wK����<�������$L�&�R�]����K�"%�cf	����[F$���[��{(~�W��ET��&��2����z���}�xO:�ŭ;�K<�' ��xF� �3ޚ�4zz�n�
�p�Q�?t#��Mg��a�vi2��y�C�
i��>�]@b��7!flB  �yD�Č�r��MTV0OG��䒓FqԲ=v.�>|x�ڌf����J#�`։��l�����E�|ݪ�ƶH�zXq���j���;�~�1ٞ�����T\�gϩ(`d��x���� �ɋ�`2�H?f7aF��
Z�t����ߩ���I��6T�b��^�<��ic�b��G���-���o����$ज+����N���ʹ�4�s�O*ƚ�+쭍5T0��,�٫I	��I�d�z\�3��C���XX%|�z�O��-8�7wjZ���?�ĥ��O��=�����\�����-��o/�ֈ1�Y������z��(?}�1�@b����P{�hY�n�d�N.�jn��>I�ԟ9O��С�<�+��,;�z�g��`i,䍣&�$/�P3' Pw��>?;!����&��2m��ED�	��A���@���lR�HQ��$����P�÷uU�>
��\t "��G��NF������j��Qآ�p�[-�w|0ks�&����cj,���@.��q����k�bZ��br���1�VdD�!&�6�1������!��ƻڒ����Rt�Ny�r	>�( ��8�v��CEq���/�:G��mi�|�f�������2bae3�����i��:)8ZO�-2�}��Z�mg�r���	Bi�n���"V���pE<�Wz�B��	'���(���J���D���?��8j~VI�ʄ̕Ӣ���]�&œ��v>4.�.(�tU���=�w��?��'�E����r9> Y����=q���3�tb&蘿?�i�m,'����ǡn��C�����!�d���C_H@1~?P�O[GvE��C���J�~+�9'nR�S�� Ͳ�{�����1.ɰ����� �)����F��!U�h�g%�y;\E��Ҋ��+���:�p��w����75ڰFB��:9�L����ΫW��z�	d���]�W}*�FlG3�,,����ӏ�z<��L�5M�3����b�E�7����A��hZm��2c�� ��h*�v�����'t�f�����{��hV�9+�[���|I\WA�V�/g*C.*ُ�����3?-.�J|I�o�t�o�����W�QԷW�����v���(�8D��_��ơ�>�΍��Y�渼�O�I�E��JQ�	=�)���94�0%�|ԍg�a����"h�
��2M�I����R���,@3p�28�bz%/�̈=&E��{>�~=�������*#B�;,����>�~������S��'��/�6,���Ƀ#��*�[�4��H�=����W.��p�~�m����J.�1�3����2�(N��ג�9v�?)Lݠ�HD �����7�S`GH�E�m����Z $��1���zZz:x߾� ,�?�����W�bكj&����:����혾x�f�P2ހ��)L��=�Mr�~��g�;��F�8�g�ǉ�6�J> ������t򜋷�VZ�b
]�	��*�&�1v�[������͞}�L��XlxVHYEB    fa00     ca0�zw�����e���	s���,;2���3�sx)���#n�b�Xv���P�Cݟb��sG)�}�b�J�xҀ��)�R%4�W��mF������"+�5y��&�0�8�P���Ws���F`�����&����$�Ԋ1��C��!j�>�lhފ6$��1�\-�,�i�䒕����MMhgj�i	Y��8Y:A�.��8w�\�i ���{9[���J�^K��U=쮲]�I�n�>M� 
�|�)@�:���kA���[���L������tnF�F��TXdWڪ�/���`�g#�1�I��U�晎K���}�1S�X������a�W�?єGx���H�	$>�/۱A��a�!��1W9z��e[W7�E"��8F�Ow�\"��g�v����^"i�����!�m��P��o�(3y�;�����D���������LUW��3�m�H�[p ~�Q?�����~_���4D��6������6?Z�ǡ��;Θ�薭�}����'(��3ˢZ�����2bl�#�w�`^r�Ft�`����9�sH홦k{)���)N'�V�ߘ�i��K�������y�tl�p��9�ĭdC_�Ԡ6�7�iRۇ���Y|b�L��/��a"�:A�W�Ɛ�R�2����*3�"���R]�aN�� v� 	�꡺���
�
��oW��S�%U+≳P��1��)�x��k?h�������G9������Ϝcm	�&?�E�(20Z�n���S!�7����%Gc6c]4G�� O�v~�8���
�z�s�.�2��'
��y�_�/ ۤfz�-���X�8`� ��a����J<X��]ǚ)C����WtvT[��@i�Ȋ^8�"`�o]�}�,G�$���*9�V�Xq#s�h��ch��\������J��:��p��V�	~E��x�+��sH�85������N��)�̫H!�;W�&�s���A6{���J��6������ИZp��k�{�Qa���Olu��n����Gd~��x���;����,ο��?#a���=%�bb�&�������JD,H�Y�(�'�^(%�H�}Ah������5n�3�� �3��R+����5x��Q=��g�b>0�@^��B۶�u��B�LzVq��=�K�}o�(�&�ւ�㔢�/eo0C�ݪ�lЅ3;����o�B�k	�e1X��ԪqW�f��C�p�s�л�B8�j���ɞtc�/��٧c��wۼ��2<�R��&���E�������ڣ������ Z��Yh������fW�C���x�k�����c%��	�&*��>�=<�Jp�]��M�o�����g�*�L�t̛���I���h��m��{<�QVYѦFπ�T��誈@AB�	`y���`������t����W��`�e$�{���r�}����"���(�Sc��D��կ�
?;Â��,��<{Ê�]!��|}�(F�	9xy�3ꂋ�#z��R� ��ⵋ�u��;-v7t�����LI�����
����;�6�E��u:������t���d���y�*���İtߙ]_W���I1<����\Qc)Ȋc�'�̥F�)�D"�܎c�)���ۛ_@�%�]�&}{���*��WM��(������-���*c�8�)�,5�[%��?0��afF�W�gK�惗!���}�L�=��Lȹa� 5�|sЂ}�CEt~��|�ȃ�xGu{}��۶;�-���yF�3{
��a���0:9�O����%��͹�=s&�z ���2��d�]�b�
�%�a1�eٕHԊc#L/��q�����3���T�IKbb�Ϲ��AnΟ�.��^m���(H\L�eTt���9�2��z�b�,���\����f"��R6n���8��z�8��� �4����C�gA�`kCk:�W�}�������e��LU�\�ͳv�`ika��_���۸�;d'�f�u6y�r��z���
#�{�#'�1`��y�W�x�C��g�/�w�$���i!���� _�7�M_8U�~&��I�	Mm�s�
�\�Fk�6�O�QQoTS�z�F�v����Rc�g>�������V�bR��]�	jzi��7�uG"�ҭٖ�f]�{U4�Î�mN�C�+=����Х�z�����\���h�e3[eC������Z�X���k�߹ʄ [��\��Y�^X}mo��6?r����W5]������]���|����Z�c��j�ۤ
#[Ń��:b�gR1?Żm�>�ŶoP|��s{@���8�[ڹMV���ޥq�~��r���G]��w��g��yW�^��½"�ˌ ��{4��3�����W>�ߡo`
Ag�j��w*�Q.J6��Is
��p��rf��k_U����?�Z�1�L�]��c�CS)�u-�9�c%n "^��pfRm�֘c}:3���\Z}��1:^�C�V=T)�;�p��y��a�I=�o�80q.���T���͓Sp�No��Gq�J�S�?�����J�Ǐ� �����a����7��7�%� �NH�9��b��}!�;Q\���læҙ�a�_O.�ffLT Y��1>�>�1q�:����8��mM�� ��E�_Z`�e�#�4�	�S��<z�w����f'}BN�X�MS�69NST)�6%:�-[������|��=��N#�ѡ�v��1Z6���&���J���;��ZÜald���WP��q�5�}��xr0,۟c�� \������wz	��P �6Qؔ;����yI�n�IDD�R"�H���#Ϸ�a���'��M��R��4��+�a� e����l>Ѯ�T����iW�)?n��>j>�n�Gާ/�&<R�����ȷ��($�Q�A׻�$z8�	���X����QS�:}������X��'U�#�>�Y�?�^�N�V�W�u�^��E05��d��ҥ|f�1�l��%��w�Y?����n,�;9�F����#09z�k� ߽�ä��H��>��
��O����	T�E��ל`������0TB��g�2�z��Тq��>*��&	r�����wT*��$����<�A盚��B����(5�&���N���)o�Óyy(�b�I�F�S0#�]�eq>�?N�j"���1:~�$�(�=�G���@<#��i�&�3�%��m>�5XlxVHYEB    fa00     3f0���_�z-";w��sݼs��=J���cy�n�g�J��t���"+je��q�xex��Ƽ# �ApZ��C�f�%�?� .��i��3�Rv+�5|%�PaXu�����vB���|�d�o��8��	���J����n����L�|��1���W���뷱~���yzf�D�`icS��.�J�w���$�ʧIɜ���fQ�RS�+X�,����S}��'�tk%e{�e>�=��29��1`�`([Om��d�H�|5��-	^��1�i�]�?��+!��!i�>l��ƋcXc_w�,�z���|��њ(��N��W=�V�J7k��O(�D��%�j�įܲQjS[���3�N�o���usa�5M��C�%~�໒Ԗr+jf��H�
���W��� t��c>�G�'�0�6�C����[���#��E��n/�ӗ�~��T�ْ���	�H��Ry6G_Cg?�H�fY�ԧ`��+����O��~�����Y���)�Ԡ��82)�>�^-Vj`�P3yG�s༨M�Ĥy��)�χ A���MߊQ��,`�K<v�����[[2=G�g҄��'VK"$���`�ܰj�e���������n	�oc�%�B�v���}*�/-?<?*���(WP�y��UJ�7�� �@�֞�i喩�X��	 \�)k򳥝>��O[$�D2�Y��z�K6<���p#����,!<�$�s(�S���cB��:E;u�=����]�J���(��g���=��)1�>�F���MA�M��Lw��D�>�q��<����
��ٍ"\�bpF<D?9D��l�4/�_p=��A�k��K�]��5p�{xN��E������b.P��ǬR�Y��|1��ѻz�������9t��9�h�{M|�YX�<WȂ�!5�%���
� }1WZ^m]mHO�N�"ܜ�j�{�-��B+�]�����dDn���O<����h�m%���q�fN��u�}XlxVHYEB    8096     b20�U��~����P@�F��R��]e���B����`�T�[0.'ޏ���s���D�n��|l���RP�꜌�O�%��;��"m��\E�v�r�zS��O��+1���&�s?Y=�?-�"
�W�}�#p�1;ܴU�k�(
w����_I_gϓS��RC�H �x;���즭bU��U�����sl���҇&|/0�Mj��z�*˚�.�:�6 ��oQ��+��i4�/��=^l����+n'��40Q��Hk�������T"������� �a�Gqa�>׭ pT�c��I�ϭ���	�@����NqBN�O��cs�u������_��r�&�Dh������֢ie�.�]��*�FR���
�@��g�⠽q8>�=mh��uX�IG�-� -�;TvrA��Zr���~f:�pߞ*e:Ia��H��]º7���A��0�@�5�����uxBh����|koב,�ᗢ���R/���y�+02��~W�~��D�T@���Sl,c�>5�o�WB�oL�n�q�̠�.8}�R��ݚ�Ӹ��%]L"�-B��]S�����:�ء��.f����Y��\����lg�
f��"W}`���|Ӻm�4�_ܑ�r#����Eh��f5v�6Ao��|W�	���PV��"O=o����?.~h^�Y����V�30(�����6�z�#�MgU�h��;;S�GD�Lm��*;�<g�|�����{�U;/Yxr��qdzQ����P?����U9��/ ES�S�N�F��t(�Z���5"��1�osN����Q�]\߅���Gn[��7Q/.|mw�x#�g�Ad�H;Y�~��z Ҭ��3�������Xh&�K�T&im�&_�B	���D �ABɑ���
%�m=��&���ᬇF�3�|%m���^�����9맍E�[d�b���0X��;�q�$ܿ�~����l��I�$���w���{�l������������0�&O�wc�������|8���� ��C��&g�l������/
��m+^�L�m~r�ᩰ�dN{pyE����G���u���0��^�����fc�Ȇ�*rVC�iޝM?����7ZkO���F�u#�A�N��V���z��~2��Ⱦ���K����P��A�:r���SRcL�8��Z)�r��|��]%�( 2[��a�5�`�b�'�'³O{�>�� 7�5xG�~��7�<	i�ic7�HU�I�qia8��:(�݇����i�śU1<��Q!k�V��m@a���D��� ��mT����c�+P���e�����Q�W5y�%��PM5R�ő���ݿ��^ߝ���'�Bq70�^��k^�ž�ce:�]3�Ǘs��pk�X�t3���O�t�F�%���ň���X\����E�ʾE�n��z49»������w4X�^p\�����sҗ:Cc��(�~����|9�~V�(C� F�87�W8�=n`��S_-���~�z�k{��o �?5&,��7�s-b�}��
*w��4�{:o����d�-T����!���oL��T)�??�\�T��8�/�-'bnO�g0��X|���Չ'����_<?\�R�y�d�!o��xߐF0�zϠ���w�_��E��Bk�[R,|��)�<�ہϡ��
�'�n�ϡ��b���0�.�s��Ȩ�Ra����Է2�z�;�5��,���m�N�N1����+��dY`i�]�+���^J�t�5\A���S�{�A����+�EO)�������n��5�67\Aw
w�L�"[�vT
��Y��;�f�"ʅ,��ٜ��p�؜:�C%]�d�1[p�ʫ�{�t����Y���az�x����Nkۉ1�l��xj�!�$����ӴOiAd��w��0���@ry�k����,�5�D�
D��]x�����؈�ӄހ�uO�6bܻ�i����~F/�d��,is��$�r(fu#N�tJZBky�Sۙ�(�{�ʸٞx��n��	P�j%z�A�wWd���M���p��nw���걄��㞋�C�F��ex�3�5���T�	� �*[��V�W�����6���O� m����a��j�*e%3�'74����QB���=_�Ͷ����Bi+�;���hǕq�CG����g��?�N7*�ڕS�I0�K�&����N���h�R�4�X���l���M5ں��1�;�8�`__�	Œ�/.F5��.�j�~�0��[���ef��ʽ�Vm�|����S�E�[U(�[�GuC��#̽�����f�xͅPSZ��W�*i���#�#^�W'�o�gM�Ui<�~ڞwqޫMㆅ�hϒ{�)l5�I������Y�����-��2#?�g0m�����С/��Q���T�#��)��2���L8Q^6~,�_�E�Va3m&gb�T�'�bo��3��/�L��n��	7A��yg
��F4��4���%���ַP J�'"
JH7�Nr�߸�U��fd�����G�Zp��Q9�O5�8O*����F�n�`�z�{�'@Я
͵ݠ���r�q0q�m�(�F�7���T*�w����8�У:�&1�98������=���>��ٺ<�1fnP��!�T��Q��.����)����KA/�/
��8���v�9>����W��3?���ѫ׶�ϥRr9�C��r�t?�A}L��_�h��!&8�TMi�8�����T^�x�Tɲ��D	���Y3��:�/n�~���à#.�މ�Zx��k�