XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����������w��AjV��j��:�ˬՈ�H�`��?x��Η/��+)!7!�Ζ�J�c�N(gXF��P��z���z�@I��?�'��e�8�p"ߖ���JKF$���s2�z&pU����$ڕ�@�q�w�.�k�t���qk���U��֘}s͍��x���a5���k�ƃ����Q{I2Z�왣B�\�I�g�;I��&��me��O\�U�',���d�sk�"�-`E�G��E��ȌS�#��X�#N���~Lk��X�-n��(����ʊ�^��A����u��-Ɔ��u��Mtь9���G�d���*���Z�o�T�e���1��Q���k����ME>~���(�)eRb�[�$�ktY��X7K��Z�LF��M�t��.��O�n*o̽��N���a��#����L��ʛ�͸���P���T���\e���a�9�swڂ�D^�*�y��;b_)
�Ό��S�+��
��g�ZY�.��+s9q�д0>\����*Cb��Nw������CB��I��z�ʟ��3�q,Z$�CEڙ9ۻ��Ra;�����|(�*���;X��k���~�)��r0�����Rf��UO<��#��7�C�&gJ'^�4 @���=a5���C�-�~�EH�J�Z=�G3z��9�D��3,�(�Հ���Ȯ����>��_��}MzB8��$S(��A	�?�� ��D1�¼��n�'���֍��k*2�ch�0=a[��9��rӖ�J���/���	ד�XlxVHYEB    5e2b    1530"��(���qP�e�\*r��TE�Ɵѻ�\�h�x��3hB	ia$m��c�i�YֳO��SR�Ҙ=N�s�b�`�#��.{Э7GH�Z��.�WUx(y�}�F/�V�?�dK;p���8�#��Ց�)�j̡Z���G8�\� ��1Ԝ�ٟ��:/Z,U����c�Ћ�O;��6:��/e
�)dR,�F�p�bݩ�|	pøy�ͪd�q�E���bv�c(T��/5����Ύ+������ޚ.^T4�Y��D�$�|FE%���F2�rm��Sn6r����D����vU7�=�Gx	�UaI�(�4�\ޕ�I/	��[�n}K���_J(�H�8�;3�d��W��.&n
l��9��=o�%{x��`�H�BX�����v�d�%v����'nEd�����3��P�E,ӏ�[����}	��!Р'�=HѴQT�g,� ���rI�&�\��s���2_�&� ��ұ�fm��Ǐƿ� ��6�a��?U����9�;�+j��6����B^�fD�y��HU�<3a}�HCܨ�ȋ;��6�6���fmڐ-�ڠ�PH�6q���ͬ:
z
����n���3ܝA5��W�=?A0����q���e^を�]7�LriN�.-X����S�js6��S�a���� $R�7I�T�z8̎����8����v�v���1Q�����=@]>��w~^��/���ON�B��~E�s��	�V鸏S���RrԮ|xQ�?}j��/Ї��h�'Ӥ�~��~\��3̜
�vEѡ;����<��x�c��Hb�D]Ù����!�J�Pi���׻���\X�r�pޕͽl�vR�U�thf�Q\|����p4׿P�K'�"[yp[��}��yEքMB(�S��fX��	�?\��ȼ3��1�J%?�XQC}��d��5�:�U�b@�fM������P0�w^���� [�Ӊ� �sGc���ٻ��Nx J��5 n�6�\2D5�;��oV���/�>��{�y1vޤ�B ž�um�!+��|���@���;�y`��p*�3(6zl��ے�E]�h����)����OS*-�0�5�4I�-�T0�A� �)l� P�j��A�Q���̡ٔ�ZS_�>�^���P�?��{[Dϧ�����r}&�kSt� �
mmU�T��ʡ���dBz�l������c˝���]���L���҃��@�R-T����)V�
cʂ���S��Qp�+�����Q�ˑ��L�������2#�d,�)�IX�2�r,���� �Z��{_iCJ�vI�]9�@�U��^%�)ݕ�}fޒkdk���#>M'� ��Qz���$#��eJ��,:R��>���"�+��>M�Vx��!��=�\M���F�7����4��i��/�mM
=Η2j�L��/ߣ�`x]lf��T���&
�f���b8��9_hR�\1��7"���6���dԌ�̀�
�Yp ��|�A{V�y�sqG�Fs��u�_Cu����6���]	Eɺ�a6dF�,����Ϗ�/t0h,����c��E�^�<t�t5���cX�6M��ɰP��ҿa�pzt����Vm>,Mʏ{�]�n��uk�y$3�6��4�i�{#�����vP+���-ߏ������D��f?��9q���(��?H�}6!���i���~h���Cg6+��ʮ�9*"%A�3�~�(���D����� >��Xt���3/NoJ��a"�;"f!��*fCY�Ck�K�ܱ�����Yॻ�y�"r��g���A>9|h�� �Q��%��47��](�`�,6lˢ�y�m��s�$M_�3B�9��������+C�4�q�^/��l�(|�R�xW���Z���̋�%l03�j���K�}u�[��G�C���BO��i�7��k��4�����Cr�eO>�s����f;qE2��(�>u��m�J�ty�_Lw�H��f�5�"ހ]��q�6tͬPA@/�MU�K�;�okB?q�x�X𽩫�;�8�*�,�c���g����Tj@Jp'Ha+s�c�yV�ʴ
����,�sS'�v�{��7؉�����E4���V3z}��f�}ɻZ��du������P]A2ҨǨ^�v{��yX�NL�M�a����K	 b�E�I�Y�n74F]�1���W2��6#�ŎZ�j2�@�g��k��+	ȁ%��b�)U)�W(�	,a^���Z�7`nif���C��5�l�D�1]���}UMHNfƺ�]����������=�0�~0#�d�;h,��[
��Xo��&��4b��s֛�w~@�	����$ld��U���O�%?IB��5c�-1�Xϓ����?�Wt���O��ꢴ�¤����T=հH5ϢxfN%+�e#�Zt�P�ȓ�a�P���.�]�|��bP�$S`��Y$���v2���c�5��������̥?'t��5��p|.VГ�Y w�$&��L.F�\����f����O��4���ц�:�8dXX���6n��6+���RR6B�W%�l�*�V���BpX��a�9�:��o	�4?X�_��y�q�Af�J�Q^�&\�Б��R�b@w�|XܙϦ���:j�XQ�t7�g��hE����)Lg>�ʍ���Y�RyB��7�f˗i8�`��~��
z�-�Tt�RA�� ��0lq�3�IM��o���!�oEu4�� ��6���
@[4ܭ� �Vh5��{�\�<	 �-˺�a���`畢w��j��L7�»F^���۫��=!dʚ���.�<������4UC��q5�{)�7�}�q#��N��o��Q������?�MJ����q��7�4\r�J-�u�UT�J��?~�}���{�q����Rʽ�$=��o�!~N���t��V���j է�U�,S����aj;B�����5�]rR�G�p,f��c�O����ViH M�7���m���ʠ����8's+����S��u�K�����X2�`鐓}hX�\Y�ȟ������1���<�2J�.��}ּ��P3Ǹ�p�avUG�G��g� v�$9:�g��@�=�d[�˜~"gD6>\�������{ΑΓ����Wi8,���+?x���+B�I�9�%>���� ���%�s!^Ɇ�Z#��$���9'�b�ްR([�����k���ذ�Y��oS?�Za$d�\�q�D6^@�Ѐ�N(�{�YC���<ŭ�^y��M�Z��&MgG��5�gߞ��0� K+s�-+�eW"K�!1]S����G *5:���;Y\m�ͪ�qԱK1�/���f���cpfx;A�UB\�a;�ò�J���]'䵍2�
8�O���p� >N��yf���-P��k6��j�Z~���=E)������-�����l	����!�����y[͡��Ũê�	(^��f?d�}���DN���b[��'Y3Ӡ
m�l�3��Q�l$�	�s�K"������'Z��A��/`;��<�N��]� ��=��_���jJ��B;�2Z���;��`ׁv�y�'>�{}a�	�/���"����h����h�)�@��)rצN��ӇVD�,�sb8���z�� .��9�:_D�N��H�jP]������@�QU��v^�ڼiƳ���<�{83�;N������W�^���JҪfP���\|��aWPur�z��B�� �;j�g��V�dF#S���g7�˽8%Y�\�	�IOo��0�;�P��a]�$?Y�\�Gq� ��1�e�T���2De��ZQp[�3�5��G�z|���� I��w����zt8{xK�f��݇Ìm$�����E9GN�N����}��V����~̏����Nm�� 'D�gǍLM�^�5�Re��b}�J)�Ǩ 5CT�^�>���L��Yt��-s~�#��Q�%��}.� �)���r2��$+��Kﭲ2�!E���ֈ�����p��Q	Zc�{�[iP*�,�����g��J�HO���<��Rt��Fd>���(��1[.�u;3���ͼxi�n1	�kU|Ij���(6�d�f�]���<q�k��FΫ&�.��-�����f�5%x��,���>�������g���p%?ó�_�'�ƅ~����%d�, "�&<p;�w�-����Pu�)f�*�H�1�#3��Z��	�����E��I�$V`�h`�!83��i�'YoA�=3��5s���3�	@M\���¶Y��Ya2�Ĕ�Ey褢e�&�e��X?��>}�c�L�M�h�J�RB6�3�
vIZ?J\�F���fVq;��-����j%M�����"�̂J��1nЃ�lR������Ҍ�@�����!�{�F�����g�2�w�J\�#5�&D��d���fH �٩�r����/^�v����\X]�Eq�7u�,ӧR~,���v�=b��f�����y��}GǻT[x��D:��х����C)b�'c"}jJ��/Pdk�r���:�4�)�1�A��|�U�mU33���0ڶ�d��t�*���������X�`�L!�犔n��g�0�<��V֬; [0��p�Z�(&���2rwp���;ו�"��ޤiS*7�`�Z�����9�TCEx�p_����@2�RYE(\��q>�B�/���<���
sr	�b��)?��:Pv��rt��_�l!)�J������|#x K���q�Ѭ�醯3ҟ5�,���;�M��u����Y��5W$����.����F���D?����^����s8����O�ZB�X����G�L]������=Y�NX��h'Z3�j��J�'�C�л��������aO���5�OE�E��Ԙ�9����X��!���.��!�m)eM%ҽN^��t�{���_�����зQoc����z�J��#��ɥsB�b:=k�mu����(�	�n��ɰ��&�0v����q�4�+� �οW�����ghtrv����Af!jL� �[H΋*�4�r�|�'�#�'�%s_�t����a/�
���w{0���XK$�cV���3�<�[�d��9݉���s���іr3������5�]ʶx�+�^ڴ�Sb�#�v	b���1�h'P����׾gV-�9J��/t2kh�c�A���&O�0P;�\�cmͭ�fn��UK��G(}���OC��-&�X'����o��:S�umۏ�:3aD�'u�O�`2�;@�;I�[E|�2S�W��Q��ٍ�/�O��������O}�ۺ��b�"	x�&@��oM�5��m6P4,�Ѫ�K6���3LQ�������/��`�ҁq�m�e���