XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K!8�+�q9�ڧ��4�*Ă�0���jśq��H�E���Tb��x΅=�� ������$y�:%�	��] �pe��ʖ��F�^����4.�F�@�x��N-?+/�f,O�Hj��vp��S�|�����Jʃ�,�C2���M��R�%-dKֶޥ����	4����t?8Y�cΐ�A6)���/��r&�sՐ��t�E���䀧�rFߑ(�WBϼX����������)w����o�jǝ=<*hWj�9+�g��u[�E����ǟ��i4�Z=�HYm���l3��E��
��`4�u��p�c09�}d��i��x��\�8�E�O�
�����͛ĢG�Y>�����6:��A�o%Q'SlYA�(�LXG�A�>�&�RP`QvO0*���n��-ω��-4qu��֎rj§�:�R�~���j۷v|�<t��Vao�i��Ez΅�
��$�ii�ŭ���*��	�lۙB������ܤ�з�����/�1`'4&s���X2���a"J���'�h�����^T�Ica��*\��v]�dXI%`21�h�}}(6��T�t��dU���ܱ��5��c3�0%�S���GW��极臠�h�?�f�w�!]����|~���o8���Vla��X���QO�Q]L˃�V��@�c���
C���;�M����4?��LH�f�t.Z��G��j=��\�FZ���\�e�L��y/BZroV��"6�kЗ���[�W���:�	�Mv�#�XlxVHYEB    70a6     b90��0y4-��W�%�1�{0��@�n���tŖ͋Y@�_�)�=���%P|2�\*Ҟ�����;P��Ҏ����39���W�nȏa��:bZ������8��'Po�'6��$��/�}[� hg�)	xp�6��w������5<�I�{^��ב�N�׼"��,���t����1'e�q*�� "2�$�Q�D��R�6~+q���}�dF������or�Og�-����CAd�)��D�z膵���оjH��@ �u�4X��x(���Xx��{�����p;�h2�x�uȫ�3�yH��(Z�P�� �@������������s^��>�f0ھ[�4���4������Ia� �⛼����m]}�XDh'����`�	@'W�{׶��]s͑:1z�"��U�]xP��V��E����<UR	������OBl)��cX��������|��<$|�7'�%�Ù�l۶h�?���Jxx1�'���X-���@ʺ�ŧd�����S��V�~#�n��u&��*t��ơ����-i�Xh��	����ʘ�֋��7���E���ДA�;C�F;Y���0����]����"��{>������Sa�S.J\Z�r�����)����]*̓��@bX�>��c��5ƴ�ĸ�ec�l	�x8Ƌ�w�O�32���o_,�����.j헌��v��	����=��w�T1/�ʢ����Q/��S5|���B�He�-��Zr���
�0�^)�!�[ғbU��&wh�%lG�|�ڎJff�=�� CA'��QJ
ܔ��[��5�b��>�q~���8b����1���TbU0���6���Uc{_3ގ�꫖��X�i�o��L5�:bH*T}��7�ÿ��'N��uY�(��Z�E6N�q��k��-F��|�yOe�ς�����C�c���	`si0zqH�1�c����'���+���/xX�J���}6���*��}1g1F�m���mf�f�,$���!��uf����!�f,�P�^$�����u�r{bR�$ v�N\Lw�3b���0fjr�I��U������f � ��g1�M��6�Ĩ��):���p6I�oq<R��ъd���p���Zu{S	֕��~Ȥ��H0"�K���).�j�>�6�Q��큿B[L�I�Kb8Ef�⩲�#��TX�9���9]Q�"{6#A'G�\�뒊��l���4X�H���Hi0����k��e5U8�ͣ��?R]���#�5���&�Bݪ�ˎa_���i�½����?skd��%o$�d&e"Ǥ?i9��`���|�u!޵ܱ��
�Nj���Ɣ��}��Z-ʁ~��ù�_�g͟����E�$���5�k1D ���obr��^�zf+��b¨ƍ�L�B���'�6z�"Wy�l�*�KSG�?C���r�~����(��
�ΞړGy�Oj�֘R%j)��nH�xkÓE�s�޸��W3�;��ɝik� X�����hXd�ՙ��0^ڴ���Ѣ�u��Q��@�OSZԸ=����U������CB���a%�%��"�n(��� �Ϣ}�;�3ͺ���.��K����vk3J��yfxX�[&6����sؓo�y�r{�xLdһ�qَ��}�_�i��/�!x[��t K��|����A,o�����Fo'tXx��"�
{�G�Poݖ^��`������Aa�f}�$���F��ͣ�K"�B�IÖa�|������^��=����U���,!���F_t$-p(��D4/l)3qw1.v��ns�=�m�y�����%H�x<)�b���+*b�J�� 1+�7���&�7���I�PB1-�}}��a
���F��搜����[CJ\��QQ����IT1\'s���j�d�B�djO�^�#�1�/��wm2�p�2ٰ\T���/O�,����I�h���\�ߣ��O�f�^2�ڍӚ��|J��%�H�X���_�\W��"f�\�ky�X;��=��n��sIJ@'��V��0�H��Kx� ���xh�5W#��Y�"��`m�d�ܼJr,�t|��4�שԅ���=�>�U�z$�?m�5pZ�vk �O5�������f�C'�A 7n>G������&��p7$*��;��%d{>n\{�i�>���uu�D�v��Β3�����G�?�ב<%y�8N���Ƽ?�@�1Ѭ�Ş��O��:\mj^qp��=w�B3~�)X*���o�����P�D_uq���T���-�f�̖,/l���nԹ�gG!��	�����N^Ɩ�B���KMJ���P�w��X��?z�\~���T�Z\+)�X���GV���v�? !^z���EO�8�H�M���Mp�sH���G�͢gK����r�d��X���ش���qû�&'qaEr>�(�j��N��ٴ=&��Յ�?�ę!�f2�ߘ�݀(Z�<��,�����>�v��!�;L��H�I[��9�i�X��O9C�-���M2��Z0�!5�PjQ;����Ì��$�����u�DA���I�mE~�3=edԭ�oPpS��k9�gq��>���^�x��pg����R�F|�l�D2w]6Ԝ���|e �$�Á2dj���ri�+K�)�k�(�'���7�]�3�U���m)�ۇ�"�� ��G0_�)z��,�5�� eck���cS$�^�h[���8��E�	�!h�Z�=�q��Y�!��|�������]�I�CY�pz�)+{H��Kb �����7q�����Vd��ꆀ0�6��9�п�}^��CY��-���p'Ic��91J�=�����]���CL\k�|�Q�t�D� ]���zx�(���������a9�l��I�E�ZH��zlq��Q4����2�/�]�i�����
�#��