XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����s�`gh�u�H��D��MqH�*����=�=�����G�� F��?��ҌKf�Va��+�B�N��j!�?�;��Ӵ(3�/�|��1Q���B}�[#,tbꔎ����o��C�5)��܈�c٪�N��h*D-w���K����C�\͔��QG�D�;��H�"iu�!j��8�Ѷ����f���o/�kQ��)n��{%�����;���EjR��d�,uk��L���4|sz\ؽ&Dc�)'ڮ���EZ���B#2;j�8�Z�"�8����ۑƬ��� C˷��L�!�\�>n�uEs�$���&��.I�l�m8����aQ���G�9TR��_�;c�9)ò��ƚ(A�%o��wZ4�J판2�:̀��Z��i@���&��Z`r��b�_�0�6fލ�ٹ����A����Li���CU� ��t-�C3@z�� �Ε˶.� v�H���xQ�̽����΄����L��GZq�%y'�o����-����ǿ7'�U�Pd��0˞S���l5�8X��x�ಏ�BW��U���[-���gr)e�<R�������0�͠s�>>ߚ��[�o��.��P����n*���� �;���5�
�_�]qF����	r+b����x��Mn	D~�%�CPX\�E��䰟E}.�q��#-[���3l�sW�M�&a���2�&��I�M㴓F�m��C��6"��2�|��Bad[�<:�)1�ҍ�3��(����PVmXlxVHYEB    893b    1e30���ov�s��E�c+��S��:!,+���`��}|��;oT)�=��)��^�*�Փ�vâ,K�؄,���"�t����rsC�OgJM���_q�뛜�~��7Ba����e<�GRK1�Q���^Rh�JAâQԽfSuAjTT����WA���n���w���ײ�bl�V:��e	�+T0�K�����2��x�U6q#��;\�,E�M�#j)�Ϛ��
W�7�O������wH���Xј�_��-T1X��X4�aI�)��o� �eB�$4 HA�_Y��֥PA����=�g��M�	��|�ͱ�.���A����ǋ�� .Hj�5���m�q�U�5U0s_��]<�e�y�YS�>I����j6ٗ��'��θ��S��jT���4�
(
��c�U�4K����r+bcR�-�У����^�²D"�L�mM̪�>�$�ԕ��5pz':Ȼ�4_�*�@��o�bף ��_<'��R���+*��a7�'��홗���҄H��30�^�������e�d<�I����
2�4��/$j���1�U��2��E�sط#�m�c��EY=9�f�[a��	��,�#E=��EEf��g�̸;�Lt#I���;��d�v������lg ����� S�)�R�?uT��2�����8Ȩ���$��N�#�i���v���e`�B�+4_�K�*�%�	7oX�ӧqY:�Ɛp���x�]Bz����ݨ�lQ����X��$�/x'1�8���?4=]$��|���NxףZs�CI-(%�*�H'�)�zM��P��`����c:�a_D�a�&�7GN-	ݏ\� s�D��&�����T�1u|�`Ȟ{�vx:�yB~Z��W�i��?� /r��T�*'Z5�:9�h �z���Eȓ��i%K�Wt!���̟�,���T�d@ml3Vx11_�;D��l�~8��mI�a���� ^+�-m��1o���y�Tԡ�Fq#�q1z��w	��=��{�u������ߟ�����7�Xc�����t��
@��C��a���*���iVUo�uMܬ������/e����Zzl�fW#����]΍��κu�� �Y�P�����6��V�[%�l.[�3
c��+�Ҭͅ�*��y����K`�?�#���x).��F��A�OŇ׭ri�
6��������i� 28�
</Qs>�^���(�M�âv`��:�ct��4
1�\WEڐ^� ���'6n�6�zW�Z�VJ�@��*H��ϐp�NJ� �R8�M_�� ���{�-��pG�;�w��=}�0I��g@��{��#<Q��nh(�g�缊��������������1��x�)u��T�l�Њ�@��~��|"�{
z*�����luj/��y��QbD�1P�`�&����䃔��D�-�}߇� �~T{��Ukt+��k7�1l�׏͚y�U��x�p��J�\]��9��)������ �@��ڠ�ۿ����d�v�y�`�*2��9���(H����iX���5����Q!;Q��![G�B��L�� 7���oϓ�hR?���J�[�/���*� �S�S�;��
Q������:�1���(�h�R��½��z�%N�#��s���`D���J�n�@&�&�^��f�)駗��Mf�����wMr",Y���#6��b���4��l p��o�|,��]K#��h59�{{Q�cj� �cR��v9�b�ﱍߝ����5�&�J������ԈZ����3�[Hm#
4��Kl�
̧Љ4>Хw�p����'�T�i��:��N(��w=[�ؙD�)���FBJ�`�F�17�T+�?aँ|R;�t#�9br@�x��?`t�Jj�I�7�B�Hڅ@�t��@�i0���@���IBˡ�T�DK>^�=4m�C`�kV�W�����"�edj�[��9�`��g��$b�������&6\F7 �X�g	����W��*�d��JOx�ۆ�}�C����Hl
d�f �w��?�j�p|��D�#Ի�}��[�O�-X��)���ho�5|8�nhީ��/hJ�����z
K��?m�l
X��vY�/	�Tl�r���e��.�/�JT��eM�=_P�) �{����$�qS`�0b!�=�Nx5�52��`��zí�Di�Z ����E�H��ٗJ�>�(�_(��J]���3�%8��B�/��$�y��6�E������w^�r5�M�L�P�\�W/N,���*��h8��w �qB�
�3�à������*0��/:�թ���˄қ�����Et���1=ͯ����>���̯i�Y��r1�%΀�!0�$�o�~\�8&[S�'�� ���u���e�9�-�\S\+�@�*^}A�Y"�GL�l���̱��
[�[��z���o�*�җ��}��V�`l4'*hQ�X�!!3ǥX��up����LW��k��.�����b�ҕcMy�j����8d���ؤ����i}$�!-����ׇ�ޥ�vNף}��@�����U���f�����a�5�9C��3e��o�E�a�kя�Jև����/����RR��O�TG�D	U�;R��Xp[6��i�����E<^]pPش������0(M�H9���9�����v���Ʃ�w��"��	`V�
-6{_n���U���&�7o�0׍�X��u��r���2o:�&�Q���毧��+oO/���.��i��#Ep��t!��:P�y*��L�E��B�E�[g�$I����*K<����<�#:�a��qd���%�.�5��
�y	 ❡(�Oe�Ģɦ`�p��&�m<\$OB��H��r0���w�P	+���0�F���/S�d'�5$���r,�:}�?7�93���Z����i��~�x�����ȇ�c�]���m�{ۻ/�+��n�V�#�P?�>��W��O�����s���0˰;`��D*[�`$�$V�V��#q(�!��=	�]�b���O�_�ؕBn���Q����ކn���@��\�{V9��T�#� #��b:���������C�ϟ�]�[g(~c��v���g����^�Z68�RRo2*Zǧ��Oؼ3�h�3�O�.�?����G��֬��p���;P��]{`��W�&�}�<4��?ܳ�3��s�EvԪ�6~�vei'�«\�;�<a��hhk�J�=Զ�z�&H�Y���=R�t����ȶ��6.��|�5v����54�i�>�)�E2Fc��24��Ox><T��2-v��Aۏ��|-��"��O�=:�?���+%�}IMe���<�w$�&df�!a������8����t�K��T=)�%�p1����O�H9'�nN�h&��@\�ؤ���Z(��ֿPG�s�-P�v�|���W���!���M���k� K#J��[��u:�x���|�4��X�.�����͚W<g�?Ӭl�A����}W[����`x5T��J� �Z��V�x�)���s�j'6�5R~�ۛO�+��mB�JK��]<��lS���w+!O����lz�r�M5U�)'B3�a ���uPF+�?5���3�M@I� ޖ��N��hvP�㦖&����N�r��8�U ��U�u�q���1���n���
�d��mx#Ϭ/�\&�T*��(p1�<������Uh���=^����E�A�y�>��}\����Ed{����ϋ�7�L �*����$��DZvw"	רU���Z8B�@�h��Ag9�!�9 Is�E�l��hTF?��K�hrq����q�Ť�X)[t�NǊw���ΡR2�?7$�L�k�|{*k(�m���{?⭎�i䩢K\��=�� o� Z�+��yT�ؗ@)<��x!�%��Qn$����`�4W���Z�1p���'3 XK ����X���A!ˌm�����O>���"s�"
ؑ����3-�"�����hF(��#ݾ�{�A+V��ԓ�wJ����V�SI\�����%�Ap~tF����r9�w��J��ge؂�	5H�D��ھ�u�W��}t�S/�����:��&CQE
O��PYn�(����i��@�������eJ>h��[����.�Vdn�Ě�P���H\�����FYgC���k�^�M`T���8q���~J�LV�}��}[��.O$�d̢��\PZ���Ŧ��Q�������d�c����E�lr	m���V[,�g�C$��ZP3��		��p֍A���X�ydf��~s���f���U�LSȭX�g�q9��|�)X��b�1q`�S%�T���0�܀��yzʿ���л��ظs|c�̘*#�RR�.���}��J�z�Ԓ�� أ�ޫ��b�(��$?��*8
�kV�I��8ej�4y�z���%v�����d��3���"K�}��3t;CӚ�l�5�گ׏ׁ@�m��I�eD������:*'μ&v�TS�����e8ȻcK
o��e�?��F��x���2�KylѠ��i=]6U��~Mz��|�`�!��Q��l���<Z��F��"�A�;��35�uZ���i��]7�aʴƯ�q�>��:������[^�i�dxo�eQ��?���c�Kc�]ؑ\@C�|����@���v�_Δrz�/`�/5�N�g.�o��6�V.rN�'bL���"pQ#T&��3r�d0_q����s�3یMSY�&]o���k�����joט����x˰i&��pZ�@�G�]D:�IȔ��׏�CŮ���Z8�=t��9�*��4n����aV+]z<rF�b8ei����A
D�c��Z�k��8`�<*n�f>��k������ ׺���(��6�-�?~�`��"�T� ����F���z�����E2�,���M���j�Q���2����o���񤰱1�xN��Yy���^�"�sk5�\@w�C��V���K��dd&��E�n��S[�p�1hu��	��38k+�����I=�-%���~��������y��+	rJ���o��n��IV�w]� �ډ��a�D���"w8i�*^����F�ԟ �D#[�k�\f���/IC�L�Ks�[M�Z�19ѳ�M����v�~�L�[����������i�(�HiB�
nyWNqܵ7@B����Ԅ��;�* l��̭Ԏ��ϫ#�iө|u$�ٖ���Y�ŝ��Ab��.O�lI��ZDo�\c��`�w���w��ػ;c���Ԛ9�7���#���>�1���]��OB �X�睉����!����CԨo���b|iD�3��x��y�2�'��9���׼7_IK>��=ɪb�˼�U�9����6u�u����*�'v�?^P3�P�@�5H_.�򐏶W:�[;m���H�Qz(�x�]���TУ'�CClR)�YA}��4}\�M� �\'����d��Ip>��N�F�X���=����V�H�;H��U�O^�y��(��@iۄ�*�T�<�|�4���X���zm��ȣ2�;4���s[��������}Ͼ��u�Ԥr
r��ԶC>��������d�~p,iz:�.�[i���4!�pr`�����f^U1\Ԩ�E�����x[�ދ�o�I@�LN鷊FO�O�}��7����K$m�6}e�u��W�������Mչ��]G�� a6�i����23LhM�9�ɶ��\���y\I�,..��W����:g\����V�����Vhu��0����,� ѶNm�D�����Xg�K�ȝY��� � \e_��Z���C����'�WN�8^l��"��%��{�R�y��2WWI;��I��Y�6==M�c�RLȍJ-�#��k�����Z���7kk�-њ����{^ ��''�[���Y�l����f����$�φ��<v�KsN�;� �b
�Q���y_(�;<
2]Dl����>�)m��6n�i�Q��=S����8�xE��`$wä4�;C�5+5#�{3
�ё����jT��`#y��zV�4�TK�%��cl/L_��Ȳa���F�W�5
*�lb���'�R�0����D��=��L��>��V�.��� ����N �����Nڲiɼ�K?qr�Q8��'��0�0������'zTJ4�0�lAZH����uH#|ݍ���������wdp�R,o+J��*��%��G$<>��Y+�;G4G=P��I��͡O���m�iR����� �t�n�'���C��_�\�s�c�1I�i�0=#�7��؅���u+��@hpP j��/H���R�|'L��s&�N���=�!�����:[�P�=AF�YMBڽ��Nfg�!v|k�ʓ�����]��`g�d&k�c�#�zq����U��oa���*Y�x�WB�b�.�)��ɢJ9��@�M�q�L�� bY#S�q��ڇ�W���R��6J:Urw?�����cu^͹L���ܗ�4��"�|�D\z̨�	�)Z��������^t��̜^}�_����L�]�;
�MC���;�DG��р�b���aa��Y�q�xZ�W����^���'
K���qf��!p��`t5.ֵO��~�+��o`�5U���f�h��=��@^cU9E�/&��_�@�	qP|_�V��Ls��X�}�&/W�]T��jv�(]��w��z��;��c��p]�i��*�蛤f49���Z�vI)DSH:��g��h�k)����	HS4��Vƴ�����b]!�����c��N��Au-�|�յ�4dk�},�@�(�Gή^�Ȳ�ֺ=���g���#��I�˶��85+��@�%�7LA�z��l�f���$<�˞P!�"�皘EFAv��{��}I@E�;�JgVB�3�'���u6��VfKk�|�'�;�K)	w���d��\��>��k4��� �(�Q��ێ�ZA��1t�ϩF�[14�˨�ͨ�]c�.Y�q�iZ���.�-�ǮaA)�:����o#7褓Pƾ� �.��e�a��6��ae8����!nv�z��qU����C�(���Ѭ� ��"L��䍋�%���F��l%���w���H��)�����=0��a��:u���G:|�ZՑ�}p( ����(3�j��A���t�f������� �s||OE�<L��\��"bl���ЄszLw}�Q.���!ر��˩��&a�oq^j3��kƩ�����c9��㨬6>�^RP������#πz��kg=�����~+��� �LO>�H4�Ⱦ!eQG�\�fO��c�Ȩ	�
]�)6qh�m��N$F4����6w�����[��em���o�p���t�[�P��� �˝�d)�ȓg^U��{,R!�Ci�_]޽���k.vFV�h�
�<G�Cϩ$=��V�˜UN�*ȲwW>�3zQW��]��HF���w�˔fO�zY?�YsŜ���g�ɱ�&�%ƣQSN2Z����$L�ŉ�Ԟ0,Zm��-��`D��-�a��e�i�5S���x�O"Qf	M�]�K�����y? 	QŢy��ƙ����Vm�f��K�lz<C�ɺ�n�ǲ+��@J �f܋���#>Ӏ#p_�w+��>��p�'R��oI�.k%=�lx\�u�v=�/F:�6�y�