XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���jF�T<G<N���������%n�J���D3sҼ�]�?�	-'o�3�#���p',d�:�~
��rD߾�3�2 R��>N!+ن4#�p������P(�C[��z7��3��
ɉ-͗ڼ�r�K䳵E��z���1dT�4�}�!��)� ܠ�)�T$���kpF/����+�4�����v�P;�H3h	�ϵH��;�8]�^��H.um��Qءc	�H��q���A�%�m8�G��[5�;�����#�i�Ev���:;��M�]��
^�������oRC�݆9�c��x%�����jUs֑���o�K� �]r�qo�պ�S#G���TE�DY|��p(�k��hz7Y*��$F����mG��:qY\:d�Ӟs����h[2������3A�3�,>����f��� ��A����2���zճ��3�Ҡ���������Q�M�2|��CHVT�{C�q��z^{������4w���hn�tk��>m;2�
���7m��$�v�DQ���"X�z �-��g���p�+�b�� ס�/o��KȚU� �N7U*�p#�:�z�����F��rs��凤���s��VkdgD��=R/4�5�s��U�6�lh�N�+X=��+�O����<J��7�~\�s1^�6�E��h93F�3zR���ہ(l�eLY��*�I;E��oJ����-��q�܏c�f�IL�V�s����L�����11�_�h���gޑO[dh���>�XlxVHYEB    3b09     f80�)d��y���&�d;K�)��#>H����T �n9���}61�B�)A���ƿ��h��>�P'|<���u�N<>�+{,��[k
"tN��h�H��-�o|�����|��u��O@~꘷zy�ͯ���u]I�l�)L��*�M�ӌ��'0�Pҵ�V�ĉ����=��;m�ȼi��e5]zJj��8����7�+Ч}w��J��\5����C����Gs�W�ٱz�o��rd
,C���P��������?�ǯ�1x��E$'��4[;�y
���n�
9R[/�3g�x�;X����`okc5��3  LK5<�ԅl^�g�u�RVT�����
$O���oU+[/r��ѯXb��0E�T?���t�jۯ�6f��Ъ��0��d<����U����W��Km�Z-�p[6pu	�R�
�I�߄xI���@a#���m?�C�I�^'!�,�6:{/}�I�v��#�� �K��>&��<��u�)�/�~���^*�Q�<Y夓]cM4�E�n4=�j�.�lGE�eɕK����}k������2-����'�&�QYn����$@�P��I�/�>9,j�
(��Ҩ������Nk/4�60�E[\{5t��庘Yc$��Gsǲk�z������o~����Ba
��C�hl�l��[�\��q�����AQ����=߃>��&�Ɍ;�*ⳝ���D�\�"�Z����<��7�h��xj2�D>��6�$L��㾒�~��O�ʢ�CZ5b�.6�J�^P��
nK�x�ѐ�]M7�C�d�u�L�SB�F=F�Pc�T)�h�:E���W2��`S��ܴ�~�fe��ʕ���p�Y�Z�I��j����G����T��%��
z�����(VĂ��^ONr�>0�;Hׁ*��Q9�����8P��\����w.�<`�D�1[H���J��m�>h�(u\�����c4��^7�����8���t����*�z��K���4����|_z& �k<[
�w�禆I��Ť$[f�
��e]�K@���Y�����A��<w�럠� E���J!2�l˱X�oT�TpM��|2�p��z��''th$��;�󔈕B��@q,�ZX���a��*�[Ku�c�G�m�+~����vsɰ�f���b~T%��]s8T	����	��Q�;�,[��v�Ń�G�O�Y�E�l4��\���<�%[o�k|X���~���� ƨ�.��6�hel�a���@�|�'��,�eu��\�n�� �(��8�=FN1��ڀ�6��\��v��Fv.����Ey ���|�����0�!q3�ԋ��y�\h��k���?B˯M�u!A/�߼w������2�+�^o慣��~��B��uU�e��fcI
�{8eX��%դ�JQG*��L@�9z�M�nz�g���Q6�·�Q��	<9Z���jR'*�"�w��v(�"���r_ֺؤ�`G��&��c\(]�f�̘w���@{iS��<�f�b,�m���4���Ӊ��l�ZEб�Gl���W�8Uz=�tЊ��,�SH�I����ξ�ϙ��YV��s�?�'���eG=����?��ϟ���$m�"�#�7e]���X��͏Rʒ���|6Ɓ��ݭ�H����XX�#��֓2g���P�ӣ�W��*�2�N��Z�s���
��9m.��Ie�  �;%[�2�j�,�I�~�PLt�Kv�j��D�����\|cz�` fW?���	i��p�j�:V���D��27��5yp�fRu�5{6�M��ej��Jn��yk�tt��I��C��@V�hP(S��F �θ�tON�|�Q֘`۴ �-�ОD�K��B�
�����ߓv�*��(-I;�� �	�[(�����Cv�A~�|,�&��6N����Rk�Ck�.��>6�x���-f��+L�u٢I���2lAzX���9|a�l~/�Di纖6��JU�Xz��ڎo��!��������7�,7���cPu�%	Z��w'��o�tVB��.&W9�:7��=S�NV��w���6��(������nk}͖��P�E��QtDyo�+F�t�g�C/����T�#���L��?O�"��n��J�i��<��aw��~�B�D�f78���NVl��~�K�3i%L'�sN�� �! �S#�`�����M���	_�3�8&�@���r]}y�׊WĜ@RT�>7O]��y؜��ɍ�B�o�#,�пP���
��} = ���{�׈�`��sQ81�n��>Oއ��~@�e�uѹi;�<�\c��͆R @��m���{û���ipN��os���D��+�r�*4�*������{~���J%Z���+�8Yhn*�N�&�G8�4�w�@���|v����oC�2Bx4N�wk�����V��ry�i|L  3���W~@�`�k%\2Nfȫ[��a�R�F5���/mf�'�
678�����*��ޟ��k� ��֨~/0�)��K�?t*J3F��d�.��hR���2���-]�0�+�?Q(�������b���V��������oo����j������Q>�l����儐d�=ί��R�Re��p�~�� 6��U����F*��� ���C=ȁ�$����i�X}�I�`7o�5�@�eIB���^� ���+����B&�f-��w����Ƚy_6q_��7ꍃ�lr�l�˥���3��R��A��^1ì����F4�o�m������~3=v���mO��2M��%OQi����D*��E-{��#�%�[yӣZ���<#"^7���)<�y۫YV bb�n���f��؃Qm��&Mò��*HOt�%�'SflRg� ����!��c�'�u	CO�����3#iz=_ ��zG�DH�ٌ�HB�W�Ab��r�X��uR��{�Q����������L�d<Ǚ�����$n�<l�]����dUh3�g`�5r�$i����
<q�n�SIdpng������7�\:�<����Lm���$��C��Ӆ?��ǝv�3��Vۙ�T�d��3�R̘�d�z"����s7�����1���fą�S�����B�O}�k7k�,1�;�ƥд�vcxc��S�S���#��O#[��?���eܟ(������`x�CٛDWv�b1�B6"���e�!���WD 5��+���Ӵ���Kfd(��c�B�s�EUD�#M@"��0�bUr�}#H|_vo�uE�sR�ʎ��-�$߱���:$��Aƀ̃/S��A9�}�D�@�{
�����F�b,DT�a 2���e�6��j}
��)�[<�K^!K;�\�*���Wĺ*�*1�8C!���?3�6�r}���Lop���K
��#��y7�>[(���ܿ�R�� �b�#jO�� Uo�,��SSX~�C��.@U{��Z�� K��XV--�e(�^��v��IR(b����� �owt���?��x���Z��w,d��^XFf�]i@�	U�����M���K�ٙ�7�":�|Yú\=���h�yb���LV�����
�^H�q��Eo	�s��0GR�o�T�^';:��m�+����>��6����&��c`�x�Խ��t90��a�A��N�j��'Z/?�Ǽ>k�y|�Ζ��5u~喡�7����ǹ'��p�!1J2'��d;�R�6�}3B(v���f�T���y��,w�5�$�Y#�F��a����E�j�Asd%v�Rukq�v%e1�����p����bNє7VS�H�n�BK���yv����mw���:���+׺��AkA6[�� w��@��ɀ�K��H�������6���7�h/|�5�P�i�B�����E��5�Z�W�*�h�0X
Mfb�/�LV�~�7���j�d��)N