XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�Q���A�5j��4: ������=CıAȢʾ�N��n>c4Sc�f8����IOW�:P�>7���[^���p�b��l��9S�Ǆ]�e�lt��1걺/0Ԍ�67���TLx�= �/��X磕J�qO��^E{� L��
M?����ꐻ��:����%b��,�i�tp7���_�r$ǐ.-�o���I_�
�P����Q�H���^sc�)���Ewp"�햚��Un~p�d��Z� uy�"iBn���l�K"Q��"I��"���0Q������1Pħ�� R+�t2�H�l�,��Z�Nz��$O]M����e2Zj7��mr�U֐���5N5)uE�%���3y���+��,"�{qr�{�)u��"�~`=;9����A���7����X�y�����Nj$�:~̟q4"� H��d.��uN�>����^�U�8	�2���o���	���px7�2�EΘ���?ld�[�ʀyY����$�V�L��ڼ�G}�*��59�$	��֕���ȑ�y�3��k�B ���է�7���(]Z41D�K;o�M�(=C���,m�j��d��p7��Mҁ��F��G�"nv�Z��a�;��yĎǈ(�����(���PXH9�KU��;��f�դF��<C.��H�t�h���X=�
~��p\D<�Qg�
f0�j	nr�{d�x��:e�d������w��������,
�d/�i�m/��-�9]���	H�_��)Vq#k�XlxVHYEB    af58    1ac0�"m��"�0��(;N����&G�iqP�=�q��Gn�LW��%� �/�#��Q r��T�w��s�h<R�v��c�[d��@�|�RI�v)�B�1`5��)�R�z�hn�z%�5����B��Ƚ~�qO�� �!Q"�z��l>t���)�l��K��H�ht|vc.��_Z}�/7.~,hB(��h*�T�ei�;�I�F41�\�ub�3+6�Tv
�#�+��S������q��{��1V�{B�5ܢ�2� �=1Ű�s�Df���S�̟�ZޮRj ��އiDD<@6��+lL�[����~r�\a4����`�ꓕ#�p�ʸ�U�D�ɵ8TB	rWS�)Y�,@�%>ԡ;�O�س;��)�U������i����nw�Ӝ>��T�E�z�MdNٌE�ަ�8���73 �X��mR���UNϴ���7��v\A`��s��Tm�pw�^�I��_�XL��v2L\���`�it�Bj)��;�I�/h^p4�����h^�#z��!�,��\ͿF��A�+u����l�+UIM6RY
���踰�Ⴇ�����7k=���q7��|��%��Xd��ugí���6Ip�X���u}�9^B�Qw��&�ԕ�g���5���|4�	��06�i�Ta�xa���M���0/-e�2��3S��(y�`�")ga+\k>^�"�a��7��jǆxX���@�dd;��?�;p��- �I	��dx��z�-0�8��Gn�d�8�q�x0���9��Yd�,uq���5� m"���"�� xJW��U5�h��PP���Ϥ9Q��G�	�ǅ�H�~Tx�*$k�L���� "�Qb���#�����>]�<m����Q_ �?`����,���PR�Tc�R���}*OKRZT_�%#�rdS/k�<����jy���5�ǹ��`��wu�ij��$�?ީ�{�e��Di�|�>!y��س��0����9]o�	"m�aQ�-D�jS?�a��e������L�n�u�"�#c���O-}wD����>���s�S?�e��b䢺�	�Nk�u��l\���W̫ktD���A.VX�ȗ3�����wgyW�Mz���G
��,���pf�2�00����q�	�s>��mV'���J]G���W=��[Q��m����R�w�������������[�@鍵�vK�`(T<��@e���R��[����1�ҭM��1{��)�X���WE%�)d�K�S4��g0���%���"��\�.�5�G�H����rsWȭZ����51���Q��(����'�Ǎ��l��nW�%�3���Z���J�N��&z�i���/q��&���^Y�f�C���b2�Uu� l���T��3#���{�d�����\�WR��Q,QL-��p�	"�a��M�+g�H�n���w��\ǎ��W�^�&7��n�)D��U�
 8k�O���ԏ+n�S����Z;�@���2�'71
2�iV���M�c���ŷg��Iu�C+�L/^'��l�u���s�����q�ZP��q�.�;j��6X�V�H��M�v�KQ��C��;��{W1�_�7��*�?A.����uf�&�gz	y���.~D�p����~�DV�@����; ��~#�Y@����+.�����Ä�M����`o/Z5�*_�D�#e�KÃc^��ug���#T�Wh��&�2a�� ��.��u�-V��X��w�و����a$P���?��8���?���c��4��3�I�����٦M7v����R$�Y)w9�697���ka=�����_�r����1g�܎���
E~1��vz���P@�Ǥ��o������ot ��>�!b�W��vm!���CPFW��~�فW$S>I�䦥��.��S'��
�'4"��l��K 4���NP6n��w�s�Ջ㣒f%�`�~+�.[jj�;��HС%PW9��h_Zr	�!���Q���	�_E���Z=�k���v�X�BS�IF��α�4�@j8R�Jg[�I6r�={Ρ�__p	=9�q確���O�2�T�Ud���"�sj42�\�t`]M/�Ӽv�bT�'�MU'���k,y����'�W��+����~W! �\��U����%�p":��q�՛��u�2�+�h=+cb݂
���M�p3��զ�^��l�#�QZ�4=����3���Fr%I���W��Z9+��bt�m�m��Q}S*@�!I �-8� �*�1��A�'l����#�fs"����ɐ��t'q)�3r'1jۙr���@Ŀ����z�n>+G��pƛg�r�Ò��^����@H��@+��%k�c;\=k(��p���{ҷY�[vQ��\��m��8�>-��P��"��Z:ڬ}w3�:��4�����U�ѵ�5�|`�ӂ��v��
����c�n�e"9��mi#�0�ְ�(F����8�[����r������Iƚ�I�����f��W +��(=*q�p�H	q��K4E�jw����o�z��#��4[��՘�.���Կ�+=W4���/�IOV���4�������qJ{,=g�f�.z��'5Z*�!�Z��*��2��6�ZWh�$�/�mt�B��v2fPr�^�j�}9�m��N�t���1ZIc�N�2��:�/`�N&6��H���:���h�R���h �<��F�U�'<��;T��7XP/��O�V�L$�cD�{�JV<�H ���`�+���_�����鯀��%V���<'���FC���U�)���sZ�C��'i�j�n[�sW�}J<���r����G���=∸�{�s8��-qXި+���������]�L�z�r��b2��'�#�Le��X1X����$���Es����z���il�yh���b:o�-�AAFr'���qs4�Si���1���ykb��q	{�Y4m<�t�DTd���� ���`,�6hX�����R4כ��!�($k��
@�[�Hɒ#3Շlɛ ���1��$�S=Mѽ$P�i��gR����IJ�L��-����;m��6�����6����15�m�j�?��-��K����KKZ�C���Z�	���\ȗ��QF{n���`�.��c�"���ͭs��Lw�V�7D�7��j? ��K�_�\��O���E���&&��l�L�]$*�e-�]O���O[�
Yt�YǿADB�<���9*�h�����j~� =M/Z��ds���W���b����^V����$ C�rs�8�J�n���RL�v�Y�d(�E|�߽�5�P�'Z���J{WLu����"��hO����u]p�ue�/��z3���^Z������FS&p�,�3'�kJ�˭��m����֓)j�a�^D��Q��\����d2���"Yt��~�!�x̯����t�飮E���xG��攐0-G�p�K�ą+6S�G�����������.M� nд	/M:�����ᄁj]9�^
Ӻ��b��#�}0���Ĺ3-L�_��S��v�m|���O�%�@�9�A�߈8�q�q�Az���ni�����UΡXy�i`X+�ޒq&P$��oa(��U�"_3Gٲ�%��8k��/�K�-�b�ˢ�k���+#
�0���u/�_�I�#߼��3�,�C\x��65�Oq�g�k,͏h�_�zKTK9g	���Ge�7	��?Ȍ��Z0�V�l�jYt4hU�*�������f�g�P��n���/���'���8���kx�vs���5j-��#�3{�N��yfY���N�t���o���������u�qp��k�	�0�)��N͖,���sa���M�F�m���ka���la��	lj����N�k��&�p�h�U�c�j�h!��W���s�{�h����)��J籾-�q����q�q�.�Z��G�Ӹ�U�V�y�^ԝЁ,Ճ��ե�_�E��_GX���Z_�z���N%���k�}�GC5|H˘�`z;�*������CF�)�=�K�ȞP�:�IP:���ù��B��}q{�c#~	�:��,�Mm[(���h�܊N�ؔ��b�|7;������t�:����9a'T�Ջ���������Z�­i��2��x��Zj���E�[(1��1bMlA���-.IA�e�/��P�,S����Yb�lAQ|آ�-Md������dg�\c�x����j�^4���[փ�$I�:�mU�Zr򞺐%�h�}�5<!"�����Db�F���_��`��ŸJ��6�λ���Ȍ�v����$���!ig��R���i,�Pi�p�瀜t��Qb	1	�J���`��#�{�GJ�{|��tᣖ%�������rdFr/�w�F����y���7RM��L2�+I�#�>x
M�ݓ���D����2���8�ih!��}��3zMw�=�f'�3����h�o܆��W��c�&ӹ��g�
��w"F鉤����J�h6Ϗ�,^;ʐ��!� �@0�m��l�lj;��u���9�]���wO�� (��<�,\�S@�{�HQ�<�=hGU[��xd�{L^��8��rH�y7��������()�M�
���h{���BcZ~;�F�7ʻ�~�؄-"uYk<���6�� JqFT� D4�q7��j���{m���e���W�!�4�7v�����]h���տr��Y�Ր��Qi����'�U�l�-���"[Ώ.����x#�x�5��.�ٶ�%EFJ4[V�Jah�Iz��@�H�}
�
�ᖇn���f�0Eq5pR��P����co��l2��i� �cϻ=�a�����;�v��#BǑⅯ[ꔰ��a���?�!al��D��w�~�H��Qܟ���0) 6%UY�����O�k7U`�8�鬫n�P�3d���@���su�gc�[�A������:�}�Q�ʸ�k�'E>@�h� ��#�N��:�o垮U�J��t�i�Q#�;��=��W�c�a5'H]����ԒS����&��x�@�ɖ܋l�,@Y�=P���	e�g��>f6��Z$�X4�ߌt�UL�� ~���\2���c����!���lb�Tm!pp7�t��V���	�u�p�R5睒��2�)"�<f�� ct�Q,m�l�����/u��@�;M�P"�|���ZIq��d�J�,>��3��^U�P	>t?a�A�wU�ܷ�B^ !�֓�׮��|�x4���b���v	��D���q��l�ic��R��e박�LAP�oq�(EJ����D�1)!����"�=>R�
b���Jj�����U;�����Vf�27W%rPt�uv�����tA��xx�:W�01q?=���?��ָMtL�w��8���exQB��(��4�Ɖ��#�K��"Q��'�I�ٳ)�e��&�q�(nz���Ou�Ik�˩Z��cn��ap;Nk2�Px����� �H8P� v8�ѳ�_��ܤlm��鏵��M���eA�"�Z5,�#�������$�=F�@A<*:��Ty��� �
��L�`B�*�U��Rwi�f0j�(����V�M3�V�>.N �&~�\��g�u?Q*Y�{���s��>_	���a��v���|�z3z��o�A#2&��.;ga��x�&k�~&ֱ�]�+uq8Ѽ:n�����ؓ8�����/�N]��Ƈ�P�n�&7�t��zr�-WV�~$C���R8_�ֻ,B.YU��#�!�_���
�����q��A�=�$�B�P������G��=������%V;����h������V�����iũA�Oل`eV=��t"\�Ä�x�xq����[X6�4�?�UL�n�(�^��p���9J�H��D�F4_dz\����_��CΜ7��,vC��,���W)���t���G�N�vc+�6d���CP���i��+�;bյ����O�[���KF-�y]�ѡ$o�Af�����v������.`h�U�OӓcR[~�ܰ�Jɡ,vJ���N=���]���)ql�?�����(+�V���YB��#���0���͚I6k_�{�ъ v���/Ɩ� ��K�ueYY��@ r}N	y��oxS�������c�ڑ�i4��{/�ޯ*��lw�k`E�L)��i`}����V)[a�Ƞ��v�8AZD|qE�Hm'?$<�Rf*���w�=��)��MV�.�9�IΠ���>�J���3�Qf�g��y�"���h�*� HBH�E��i2XD�[�!����h��*0;��r�	ܳp:m���ug�4�����FM�
]�v����@��r���.��P�[�E�!y+�Ž����XW�JYE:���/�V����KSԍ��'N���!A����H2��~��\Ǎ�!	d�ۉ�MF� ���1��\ z,9�b'F���>�
��PL��O��1yE�1�qj:�L���'Ҟ/6��� ��h*ێ;F̀�Qӌ��#/9̏5=m�(�,�KLi��ً3�P�?� u�nK*Ԯ)&��4/�:��GN�%�����S���y�}v�����{���<	�{du.P9�$�� �������lzLMޗ \�D,��w�Ƨy����t�:�&��!*t�D�G�3˨ʣ�3�v��#z�>��pUF�?���u�9�qF�.�:6#�׳S��ϣ;���e��j%�V'!�0N�N��m�*�˞Bd��F�(�fH�q�V�2�ϟ���{�
m����̢P��"4�=D