XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:_{-C�h�Q�NK CÂ�>n�k^̥��J��c9�ETg�|�mu���;Tcz!���(�$�2*�����mL�b���R��E��NޕƷ���<�yș�m����뜩,�}U����H\�`,f�<�o���opFo�*��QG��=9-> ��b ���S�Ώ
8�_O����(W�o��I[��J��zҤ��䌛�b��Hlw}O %! of�&�$>����~�!�K�UY��-Z[S�QL*�9��?��5��Ce��g{���a��yZ0m���ta^x/��y-�͛=��Kx�r4>T��ʪ1`(��>O_<����6���TQ�!�jN�_�m���ܙ~���Mҫa���t@͡�~���(�j���c43�À%"�0������綯������u��9޳�(Ǒ�0���A��P����\i�m��*�iA��Y�ɑ������<����P�q`�����Z� �|��b4L?��wJ���A<�h�E]r�2��j�\�H�67�?pnU����jG���2͖���."��D�Z���}�o켙�U=M��^�wilĿ��c0xbiT��z����%g��1��v���	z���[��љ� �w����5/��؍��"����
!�;��(}�Jh��H�M�]�h�7,�I�<�A)#�Ԋ�������N�x:r�;����:�����l�7�'�g0.���U�TE��ޱ��za�J��\���%]+m�L���Is/��*XlxVHYEB    95d3    18d0%�IB$R�����?,�>Fp�f�hG}��l�m��������	kQ����g�9i��&S��B�/q�Ado��<�u��C�)�LE���4d^=�<A�1��c��T�Aw�C�BT�=s����W/6/O0TA�<1L�&��1¯5���;ȳ[!h��t6��~���s�Й��p�zj�`ÑL߽)G8=�Ϡ�۶5Q���
@x�#g�V~9�ړv�������(�<��c�?��?�w��u�u�
F2q �s�����|�xt%�<�h���������Ս(f7�}&{���q3DΟ,��m�?G,����΀`P�+�h?7[X��+s��#t�s�7�[6���� +M�_=�����&S�$��SgwFG�.`×͚� ��u���<���7��+�6Ja]�׽�΅ρփ��e{���W��*N��\Y�e�B'ԋ�������-�I�A���w]�"޼�|5ě�8�����A'�s<��c��x,��d����%��3#nۧ$+���|G����|ӄ�6��훽y��H��^��&��z�騲��i|d���>E���R�T?_Q���9Q�X��Ԡ���W��z������l�˅|Q�����Q�j��|��,(fI��Tp��C	���t^���f&=�@
��|9��oq?O����[W�zDs�O�U�o[�q�8T��.=��.�,����:�A;���dk|FH�����.��$Ju+����S�/��ѧ���yH?��K& �Y^���^n��޺p����*��[-�%C��wv��~�)P���d��is�^ڇ����	6el�t��C�v5����C�P���ŔB��4uf�1�dHŢ��1
�pBJ���n�Ŏ��lK��RN�'�"d���W���l�p�~p�
0���vƭܮ~��5�Y伅5��M�F�N�u��^ŤǄ{�",��VI}HA���j�O�K����ǒ����]O���(�	՜/�6fÞU��?�{^l��<Ђ��������<N��Z�J�f���-�@H�;���T�]�6|ᓲ*�:wL"�㐥lɭZ�"$Z��l ��snQW�&���,�B$2�y��ᙕ��U�*�չ�$���w���_�ͨ?�+��PB�ӊ���z;Vd	�"h}������v�E")L��H+�qӟ���3v�ֹ�h��f���~��1��X��l�O�3�`3���f�D��Utxiu������J�]۠yv�n'�8z�^u��_���!����x�ޖ�[�Qu�xy~�w��,�̉�ԟ�j���!hDngk�r9u5�sA�\晄�>�p �#�Խ�7F���>�w��~��u��<{����Ly�ms����}6������1V�B7��O��T�r�g��f�א|4���l�:�����,�la9��dv$�{��,��N�B~ÁPý[t�x����M�i��j�u��G6Ţn�x�[�E�P��:p�>���Ɛ�8Ec��@k��7���2_��pgR��S� �^��=�ʣ��^g���%��D���U�f�O��m�5E��`n/��x�Ǜ%�Ęf0�V�}ms8>dG�<�t幓�
q�1��}MxS���w!��Y�>�c4���kW�ժP��2*�6̳P@���uޕ��(�z�m������a532rdD��4WQ�0��5�;\&��ÓC�	��^%��&��j��������!�'9ڛ�B%Ց�`Y6S���ٳ(h�DUv^^� �V�b,�D,�ZV9�����ީ-��<7��:4����:��e��$ﾢVcaΑ�ej�V��9�I�ׄ��B\��Y�}.N�O���x~��y
>I#a�xϊ�u����(�q]���˽����'ȋ�=�X�4�� �Epz��CU_��l������q�>��_[�#�Q*mփ��S[��5����K�t�X"�fڢs�����-I�-��4?�7� �&����#�`iM��%����6�mN4ր0f�g� �el�ű������#��N��]ݗwn-��9�6;([�&;��x�}"��b'��HP3��b�U	�C��!���Ɣ��Ѫ��e�M����UA��S�a��ME�N��悢�`!r�eGg9��u�	�e�Pe�a��8Hҋgd#��!�\"t���8Y�{^��TM� r�x����r����w�UAy�%QP2��2^z{nmW�a��NyzD)?	#��8�kA����q��\T.��Uؓی�c��G�.�!kՄ�]�:�w�2g�G�;��*V|�P7_n���ł���ӷ�4�=���S�v�I~n"C��;��A���X~p�xL3�7^t��Z��5"sJhU����8�`q����\��0{��h[�����'�� Eӝg��4"�B�;�m����3�ӓ�]�׽�B`+�(Q^a�Y)ֵ?$��Lu�5d	�xJG�}.s������W'%e ��:Z�P3���>^4�o���q@�0r:)�?e��ٟ�l�?�B�����T�_4�MX����bá!���O�E?���r�Zu�3�3�4�=[���r�%$�Lv�yݘ��T���hp��&�K=h��٦k�8-p��DkN����RH��!���=�B�5�ң�lV���ы)&�LXC�e�r�_�Y�I�d]t�k1���7�\5��/6~O�Et���t�iV��˚�+�m֥ꤼ��c�V}W��1Q�	%�O��zƗ��c`~������H�}[Y:�"��q��Šfȼ�� �{����k���]������JE��=�Pcd�����s ll����|;n�>�"�&��]�s�ajM�9l�J�z(&��,�����u��4�Y�	H�Z�Q`E����&��Z��5(��i�BS�C&v=���~
���5�л��+��*�QV*�m�a	s�������Qw[���z���bB��>���c�}��Yk�e6���Q�ci���'�݉dt����iq���G9 ]�gH�F ��Y��jSV`�Ħå�z`l�7��r8&����f3���"��G�Zb��a
�LPg`��IC9��W;�c���lf�[y�����nSs��Ǹ���]6�����^����Ѕ�q̕9���!�<W1�W�Pܩ�n��ge�>�[#�v��)f+���8`m$�XMO�
a�)���s>1���/��-����M[�;�"Τ�����D�ԙ�����:�*��=�t��Uw���ҍrG�������� >�����U�	�a�f����`�CJ��e�h�5���e2tzj�b�N�G�LA�Yd�=J��7CG^����+��H1�L���Rp<��0�P����&_�؉~� ���=;��5͑���1�
D�֗cq9b��/�wQ�����х����<���� ������A��2g\c��N��xU�	�b�R�n��H�;�T�[�#�����1R��x�D�,��a*R	��'[?��=%⚜X�X� �� с36+1D�-o��R.�iS>{/��?��C���5-9�����$=V/r��I���]KN��ᅔ1�ru&g{#�)كj�k�
u��2�a[ނ�V�R���8�ݘ[���S��i�e�䳵��)�S��Q�=6�^<k��8���$üBǞYeX��-�@�}E�{K"xn8��DU�M<��
~&KJ�$*���������V)i�zUbw�P[~��!e��`�ƄRD� �vxV�i���  ���Nv�$5N��u������/l�\����^���*�N����[�'w*��n��}�T�1L�
e�J^�(�f�yaw�
I<^�htƕ���K2�G�$��t�ٿ�b����u�?_b�Sh��輫��h�:4�)V�҃�$k\t�8kG�V���(w�se���;�}yB9h��-�Z-Kjkr��X�t|Y.ʅ��mQ(a$35����r�bw>B��l�8���~X�p�r���3���|�-�X�(o��тx�*�<L˾׀R;� ���(����>PM��U��!�k�̫J��)�M�(��u�w
��A���Y(u��*FW_���4�w��R���R^� �-x��Z�g���ҪVx:�q�>��֙���n�-����-cѷ4}��Q�]-�V�q���O	cyF9���:��#ͻ��T�����^��<�E�}�_�����[ܒ�)r�#T�@fdh� H#I�1�G_�O��+�*G2U%) ���6�ș�wn��Z\������a�e�Or��
�
گ�/F�D"�o�8h`��-	���ʚ�S&��b��(�T�E.&��4�%bۡ��s�r_ ���g�[������nn�.�ӱ�����=�ؽ��]{��ͤ���G��ǆ�iށ�.zJ���0�bP�:�ى|��e�b��5��q���_�6Bn}�(�tN��i�+�u{�?F�襥�)��r9��k﹫4�`��@ϣ!V������F�8�L !.Z�Ib��s�l��
�M���r�����ȷ����FRN,�f���������Mpmٱ�T1e!T�?��/d�K��h
"��ۋb�-v�sWa�**��xZ�?1!�������ዩ��%1)��JG:��ƫ��dv%�Ƙ��~`�UJ��v7��#T����wkN/��.�0�����
����8�<�S�����Ǩ�TU9�or�V�<���/�	��������؈��đ>C�,7�ݍ�b��8�Q~�g$k�֠���JW�k�V���N�{K�4]N.l�6![�l%��nY�e	U�.�kqQ�=��)�@��E����iI/�qs�Ɖ{���M:|���N5x_�c��5�N�A2��$�0�&$+µ���bk��CM�;��@ڥj|rHy>v&�fS�k��b�
��?�5���-�I>3t�V#�D���#(�{� �ɉw�2SOzI}@h�6�Ϭ�6��C0cj#^�Ƞ
�Y�&N�H�p�p71s���=i�쬆���+��c�����bm1�?��Nt�ȾP1�,�h@|1Iq��M��y�r�NT'j�7d'bW[.|E�8��PW����p1�l�6��[�"2��-h-�[E;M|;C3_�"�*k��y�o�m�V��/�PTB��H�mF(*��L|h/�0�o9Of�Q�h�C}�(�����BK �3#.����L�������Ǭ�H��_A������t{E�K�0�)���Ҙ��qQ�~��r��cC9c��3>Ǎ<����w��>nÏsܙ�W�z�����[�d.9���Ѩh������8��\�F�n����+�}�b�KYV{#C�lw��\���н�p��"3\[[bd���P�k@'�� ���[�@���
SV��������F����bR���)�ft�އ$X�s�ɭ!|����Wm�B�ɛן'�k��%�<����䒤O��۫K7�{>�su����L+��',�,��3F�3|���ՋS�d���G����嵌�L�.PT���:��؊�����wЧ�M,��-![��=��A��^��4�h,��LX�E0���:����Āx��e�|��&��_��^��N�6������q$����ӞSo�ȓx5��֠I��BP&,ƮbW@�`����;�#j-5�|����ځ�j�S�/y�r�±�sⷧ��ΝV\�f�!�/1��i�r�F�nj�6cY˗�>reN\NA�92!$�C�'��u5v\��%��ϋP�:����3��
[ɏ�)�Ϻ$(R�L�W�����l9Eٌ����s��S�fl0�� @i�d��,�JIT�c-/�(:��H�;2��2��4@����E�e�§�,������}h���x��f$ @�V
�Z��@b����M>�B Aҋ����������1�?�&=���߫`xi~�$pVe�4���cܢ!�_�*���+n���L�����Ng���_�*ے���5���"\Aˏw�0ՠ�)z������%�Q�lu~QU����d�u�͟���K�@�����I�!G
�sh��/�&�;��Z�a����A��]��u�����^FL�P�Q�Z�� l���&��a��!3g1>p#��?�C��ÁL�oh�P�n4�1��o��'��(ר�GB���w�+!r�tuz:X'Vjy���6�b�2�5Չ�5����c���[kb�iҘ���}���|4FVknnڔ@�1љ���
