XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����� 	p���E�:F��`���R�Pb{Z��&�U��M��^�3�<:#ƒ6V~���zdHou6�t^j����{�N�g;eO��̏��v7l����Yjh�n�2������;���C���2��)r���D�@���"���o��E�َ�O��=	�˸����BM6~]��6Y�8&e�n���{Q�$#&�J�s���&���]L$�]����W�He�s5�^&4��W�X���tL�Gޞb3��?F��c��o����"�����Ao��/��z�q�'�E�7��
<ӻL���h��0a��G��?�Js���ᆍ=��j`�}���d�� ���UvI!т�=�`�m��~�%�S���9�p��ҫ��½���VO����Q�	Nz@�B�A�6������I��CTΓ����er������| {٠.�Ϡ�-�GiY�s�a�"���Hg�(v{~V���1�v]��!�d�[�'j/?�t��!����e�6�X�w�8S~U F�Hp�-0>JFt3������֏.�p��pk��V>OQՖ!:�lz��:�^c@�{m������e�.��X	�i˭��_��-��@�֫���SzJC!�P�˺gK]Էw;�$��z��Ί��&$D������ͫ�?G(C�ȫ#0	����)��O!l�ӏF�3"����$���y��H�nfR�!k��d�^j�-�2�4��t�٨>:$��>��	���bn<ӦB\7Ԧw�"T���?Ћ&8���3�p�-XlxVHYEB    15b2     890)	�gl�$s;@ u	"��Y$pJg0p�����~*k\)pIfU~ߍv^�£���-�i����L�o�%p\�|����6''2�Nhk4�`�b�U(�V�������!�P\y��K�կ��i�����T��K7��ܓ��5�5�Pܸ���4���cOn�T�y(��L�_�� ĶW��ߋI��A�4�F�$���ƿ���׋}�����l[���J������5f�#|EY#�_�]�3f��w���φ�1-�m����6�9Ql�a�N�U�J�,�&�~���B��������!�u6�����hp�Ra���5U^����h�O�KIYɌԌ����"$�9���}^x�y���G��=Z�0��|	�פ�4�ʰ<y}�{A�'���I_=��|������ͯ��6R�����es{�����WO�NM��K�_��g؉�i���Z��}k�nfL����<�A�cϣ�_�y���C몺%�f˧��K�Cft�6y/�6^O�,�����gegm��'��/�k���;[a�&�C�_��D�映zscҭ�0cX<�s���]�р�=|��A�ݴD�#�_����`�N1�@
�^p��VnFc�=S������0���s��q6�g�~��Bo	Y��\dO �"A%Xв���qr�4!�j���[�Q(;��J-|5���c�UO�f�]fM&������W |
B�y��١<�w���%�A�����
Ug�y
�M�_c����˂`�������Ǖ4rz"����ȭ	�d:켯P�L���M�d)��-����S� ��dUx^r.E�������M%�l�EXۀ\��Q�^7 ćɦ����������.�Nz����7��S��M	jif��HB+6V���u�u����JH㞆��f��7�=O�1�[Y�D�CP��X�>)i��`��<����_{j*?ʟ�Yf���^��"i�AJ}��ݧ�oK� :&���
Ls����G�I�OUZ�N�����K��r�[j2�Y0�X����.�����m�W؁&���K���u��Jf�#%������ћ�m��	�dX��X���3�S�:q�V�gs����q�$ [�_�"�a2wI���g\WY^/o�5��4�A7�3��m��-^���C��&Zt�AA?��/���ca�B)��|5�緮�S�E�o�?���n�-&73��֧q6� Mc��B6�L���e)~>>}��?N��o�t|���OIA������Smu&��w`
��S�9mI���-3B�{��9P���h+�W^[Lyv2P��-�,g�,�%���ZvM=@�&I> �X0gnQ.W��4�hR�"^s��=�y�t��$��&Ou� ��o���ĕ'[�Ig$��W�6Z�$7*Iv�/:v����Ou���8(T`C	q����Tb��>	rP�T�=�m򢍎���؜��z�,��i��I��G���������!��B`����h���-�"w� ������`6p��Kq�S�R�N@`lӯeP]k|aA%wt�� g"�k�)����R4Mn�0L%f�l�>p� �h�M��v�Üssa��s�YT��]�ӟRO����(B�v}�l�꛾Ik/o�;ć졎G�^\��Gt_E�jp��s��d������E��<��n �d��@B_�����O�4#E[�P81-<[|A;�p��Sg�cn����9o����~6�5���7�1�H�fH��@�Zxm*ʕ�U,�����)Ld���c�XJR�e� �s'�̧�t=:�TnI����O�_A�V4Ѩ$*�z��'2aC��2G��vv���t&�]�؟�� ��k�H#��3r�[�Eً4����]�_���T��F耪��P��ԙo�
�˔[��`��4�8�"�e��E�-��F ���C��`˭�;��L���Pd��*�dS�k��d��!P����
�q�*�=�4^Mo����H
�U�!�tgJ��>�����R��f�=�(�!� Jqˆ�P�j�E�v/3e��.��S�J�gj�7X�����Q���S��
��{��=��x�r�,��~�O��9��-p�������T*̚q�����<��*թ�r�6�#���֓�}п��z]���3{v�/Ʉ��;�Y���g�:��ɮ