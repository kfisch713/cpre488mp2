XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.^�I��-��������#������χ�-mi��u���ozIغ��=�?��vS�Y(E����0��A�s�M	���J��)ƍ?9&��q�U�.�� a\*5Ma;�s�X�HW��j,�cK�AP��i��������d,x8c`�'T�=r�nW�ԝ��v@Y�I�0����r���>N��]n.�{ SX�AV�RN�bT�����D�v��"j�.!���`���ʅw�:KT�NyIl*�_aLD�Y&-2��]#�Xۇ^���2M�%	c��4���g��5�3$�p���`O7�p������-�i���@�-�W����{h�a�\)�F*�ufUowd��6|'U=�)���'oe��{�����s{i�wN�X�C�BZry��щ�O:��M��:�>��3�jAXb���Yg� �[Us�D�
·�pN�߇1>���[���='��Vޒ�lKb����|��֧\h�)��ʢ����K�څ(`$J�	�q�$�J��A��X$ʬD����/Qp�@���B\��x�3��(@���|g�*�s�p��"*^��4C�\���BA����V�?�������NNB��,�@Z����P�@�_��5��a����W��a�E2�����Mk�R⻼2U:��#pcN�zpQP���}&JJ\�
��5�t��ė��$
����S;�.�]ˊ��GS���6�[�q�x16JrR	+�s�j��P�H:�Ů-$p,3eb���|#0�����y��[�XlxVHYEB    3fdc    1160m�� ���HK�������+�r����^�����:�� ��5ԥ�`X���&v�cZ��f4�);�'ʻ�v�<x��_���]$�|��7''��.@�Hj"b�^�R�.����!����+�����}����/�j�0os�=�/����j&�M6��3�I/:y֚������8_��j6L?�q"��� cu3�3ŵ���S�D�QP����p�[�]nlR's���LF�]=��C����څ�E���k#��GL�j\�3I�e�r�Z�,g-r���� M�?G8��KI�}�]��8!?ZYa�x0(��u; �"����ӏ��lB2)�����`��#�~�*���U�Jw��)�m��j�!�����F��T� �}&P���y@j�V�{�ᣇ2W�ǳZ�3d�l�qx.����3�9VOt�`��d��p�iQ��@1ȼ?O��B
 ^J�6-�Ԏ���uZ��X�hE�k�]��>q�Ţ�� KB�����z�r&���@�ʀ�g�������,��2v��A֕��Q��<�g5��2��D����z>g@(X*��bq��mc�f���?�����Q�|��<SrE��v��t!>e�h6��J���k�NQ��>��e�(�[�&��b%F�Ua��iy%b [��(���̤�fDh
��Y�=����#�fE����?�Ǟ������qԈK��	��;2,K����&���J�_��E�H���b�� �����p�	I�<�����EF�GQi*xe�-8
�����0r�>�I@�GU�@�Ϟ�N���:g�]O�q�r�VR��D�!��p��Z\s�fj��yG�m��Y��R��o��C4q�<q~|�� [���iT-���O��^�A�9�T�>3��y#C"�"
��(&���x�s��5e��/镾�tHq�ot��A��4�.�%��2AzE�$�p[͗�9��jC�O�A�;���3WdM��3}�:6���zo�8'4}��e~�6��9,�X�1c�)��E}CI0ᘚX����Kn��Wr��o]��*|�������h�M���qu�ϱ.��(l��3��y����<M6O07�/� }�#σZ8n��>�Y�!�� �˦���]n��bx��}����������&�j��P��S~�6Z�X1�4P }x��L^��oM�Q�Cl؅�ҽ>��-��Y|M}�1c-w!��e�6,�ԈK��(6��T�������w��7ni��;�pGDtg�����莼:�?��{3�P~�ϻ�W*7z�Qϟ�uͿ��at>]�N�	�,���K��_�;V�Y�����>���]��C`;�(pM����,&�ֳ����[U��TB\��h��E��͙�h0,��� N�]�����r�K<�~ 5!�����T��dح�&|�H��1��$ aZG���r���A
����$?veӣ`X�b�J��b�>�{s�|-_�ޟD~˘�(Kw���U��͹5���ژ��ۭ����J���B��������w⨽�G$�E켳�b|+0_n��[��#?�X�tt���􊽢��o���NE�^N��y��Í>hS��^F�Ȟ�z�����%���}>i+O��cpR��zad��g�4</_X<΢<���OJ�B�����si�@�5ɿ��P�,E�N��%����i>��a���g^�;3`p��pYS��-vz!����J�d�0H�|��/,T6���'ō��%i�
~u�l�!��q6�1�w$��3sv���!�e7�lI�|�@M�x������pUv��:)�K�B'�����o-iC�5�[�h$F��]h~�T���ռ��iF����a\�`H@��挡�c$�O�H�������E���]A̚����g",��a���:'���;�"�X�ϔv����� �(&��T�o�����Q �!k��[�. G=�%�$**``>Ѹ�>	�d�X&�׀���A>�x,_��᧵m4��a�k� h���5��.����@4�F�U�^�)�a��Bd�6�TڦV�_���2�ʆ�_�n�d�o�kk5��͛\U�@�UpE�#C����V7�'ۺٷ@y��N��P�L�V���ߨ;WWL��B��Ζ�I� �����995Q�}�1%�i�L��^���NHrߖ��yF�	f���QA�t�E�4Ww��Dƾ����a���$E(�q#q'����-�x�3�bb3.�.ҏ}L/ՕR^gI��F��>`Ր���%�)�3!~��Qo^U����1zD6Ɇb�X�t֦�4ݣ�..�r"�%���w�~:���o�V�ZߤQ�ہ|�|��Q7�r���K�<e�uY��̳Y�!���	�7�k�]��S���T>���l7�J���7�g��f6� n�'�[���at�KY��b5�T�l�F�* �PV�7~d���%18�,z���$(wTF��&�P�� �X_����'�g�W����O��I؟�F��ͻҳb3�D�Z�M�w����k�o����s���fN��8��vs�,����b���Θ#F�WXtؘd��E*�������t�]Bi)���;]d��%j{Tjd��Ɩ��3���b�I'pV�=��������Mx�.7��ʽ���O�g���~��)~])�(�~�Tё<�lM��vg(7%�[�S�)�I9�T�2���7Y���?.c�ܺ�U8\!��s/<�v������$k���4S��b3I�X�6�P\U��Z�������㾔�b�Z\'�܁{�����j��d+�����z7�We}H�� :��0�88.fG���JP{�����C�+��ֿ��o�GK�������*J�o@4��'�=���1N�s�|"��V�遍�tQ���	?��~�������S�`\)��������&�/q-�q`4F:f�.,��HW���*D1��%db᱿mV���|�\Ubi�q��ak/���	_��)����q����(Tsa�O��u��OI�!�Rt�䙥�u�7��?X���4P톒;��	�Nr�_�m�8Z�&��_@Ǒ����.6;�c��8�B�5�+��+ �(-��X�Z�`�Ix��u�au�r�M7�ů]�x,/

��>x��ǏPX�o�ڣ��<�B]E̵�j�'�*�����_B����rQ�Nr4=�̊b�rn�+rɰ�F�~���j�j��������q	�C���t��\D�1��+�Y�}��MG����P{z_�����O�BU�}U<
�aX�.Z�����?# �D�M�qhO��	���u�t!M8_ ��#�w
b$��9O��$����L��p�^�`�������g�E?�V܃5�b�P"iAlܗ��A<Ӟ`�j�<$���}#�%߶�����'aD:>�&���w[�&JZ�P��Y��{uh<c�����$�(8.��gB����ZsZb�S&�a�aYSG?�v8pvt�K$g��ߝ2��.�Lx�Hn�QN��g�$��q{�p{��2V�ٸ?���.汣�����hw�h���z6�9bF�����dɺ�5�@Ԫ9�"�D6�zS�{$Ǧh�Mo*�h	�c
� T�d8�@�����G��T���bؚY���+w��5䢝�K�\�@�,�">^#�>�7c��A�@;zȲ��Doi��b4c0�������BTQ���7��+�S��7Lf@J��O�nP������"�n�"H�XT�����2m�P64㼯���W�258�7
���q*
]��+	%�ΰo]��^!����:�z��[ՋE�BF�*CdBɭ��>��r�����b��|�7���2�;�RN��^�?�+iW�d��3��,��GӾ�҉��)B(r�fA<e��XⴋN�xdY��q�?n���y�/#�{ρ�e��5��;�6(O���:����d3**�i�
Y�U�����Ls�|w�$�7��@{u��?a��ܐ \�{�ŝ��O��{؛�QK�ʹ9K��.���sP�{�`�Dm�l7�f����˯2�ץa�{ԽJ����(k?��0�v�)m�j2�3�ц枍q/,\��&l���Ә�h�&��?Y�����H��ǂ���|���I�e�vw��@�癖)شɳ��X�����,�����X%��u��r�Ybd24�H�z�@;"�f#�|'�ws(2
�H�������t������A�eJjE!�����R�̏�^����U����V	`������,����>\��c��7��`iY�mU.�i�x�,��H��@�'���8=9<��c��RQ���G~�$��b-$�Dmq�9YT��	��KC�#%
R�yѽ���0