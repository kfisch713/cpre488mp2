XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l���eY��ȟ-�T�	I���J�(�y�$������������C��$�I�%Y���?9@f��ӏS�>�z0���{A�	K=k�!�"-����iM���w�H� �]��q-��	����3w�f�G>!�܆]�L��d����@Z!pQN�jJ���
3�*��L�-�:OsD��1j:������g��nʭB���	����y��p0O�LM0��l�q��R��m��'�����V�͞��C�px2��c�/}}��֘��\kS�
8�eş�Ѧ�m�+<����Q׻)��Z��`�J��m�&�E��"M�jq>U,�Їԡ�D09�by`eQKDF9��0Z!D�:>O!��¹��F��gꥉC��g�JHGI��щ���9���ܥH�L�l��7��<F�ܶ�����އq'����3�c{�_??�a�������B�R�N<
<������W�h:�nY$F�#g�{��^3.����4~k�f�.�����8f]~�4�ܝ����ͩ��K*X0%�OJ�:	e`r�j8�L����<������Hˬ9�Q�-W������/V�@����(������L�^��"DF|7: 0�q�����]���\��8����:�7���
V�c�`G��U������.�yl�=��P|��E3���_6�Bew�1<�j�nw��畋�H������]/0���4�ra�>�p�c��%����"+q���#;vI�^8cI�2�29:��7kp�XlxVHYEB    1e3a     a20��d#���U(!���sP�t�P4��A�?g��w�u��0����<�H�HX�q[������L�ΞAO��<sq�d;���.���A˶1ײO���G�|7��U��3'}=�`U�*�otW����RT븨R�>�J�d��O]bYͽB��,��o���/픈���$�ĵ֜N6�p�T����P�	ԩ'K�@AS�j�SK��30ͺ���]���E�S����H&����c�,mف��L�ܻ��a�T&^N ��=R�u3Ԍ��Dt h���`Xl�u��E���x�d�*p����ܳ薇~R��j���N@�r���c7��I��wL�BsX�n�P� ��e6@ߧ;����d��wے��G[Ƚ��7�������@F��t�C�qc�W?jS�T����Ձ�!j hV���0�܎�9ۿ�R�h��'��0�(E�*OAB��^�Jqh�]^}�X� �������8���J��ڼC�c��-�\+˅<Y������u��&�)���~y1:�)�7�|��a�����@"X?�����)V�0�:ل��N����_���ò��+Q�/��%Q��.[v)�����@G���\�	K����Y�����@�h�-���o#�~ῠ^����U�@�yQ�Jn�<��`�,w�t/,N��[�&P=w�6���BЉ�:!�6����9�q��M�1�{d�wK���yўi��h���@D�?�5�7�����,9�Ň��+���\�g:��țU�1	��z��6�d3褛d}O4OC����Z�£�m�2�~��
I�W�'���A���"kmۣ#3�85����"#c��-8�������ǳ�@��oq��3�K���2�=c�$<I�ls��ؒ�l�}cZKّ���?:@��ܿ%�]��v-��I �6��!��'��o�88C�Z�v���gʻ���n��|4hutX��u�Xe�3�7����&��)�({lRP���1k�-�t�ohd�tX�>ƭU��~8a�H��9lۊ�3q�Mm�F��m��~�`jY�7��F�b�;h�}�tu�y!<l^4�{V��`{��%��$��ll(�.�٣ @�d	z� �;+�� �PL
�3B1)�/{�#w��Z:��!��Ӎ/��݀�!4[J��i�z �~�k}�g���~ʰ��='�s�u�z�+��*
-�3�
%Z�N��i �w�����j�c��0�0"��D&ʰ����������K铥D��sË���^R���q����JP�e#�fYT8D��&�2�:%�"A� ���e� PZ�U�+�1:�x�'���=�BC@�5����S���=`O&6!E�[M!�nC��)�ݡa�jd&$9B��O��v����xݟ1�*/��u;@ h>�F_~zS��_�$-yk��R-�u���do�*����ìW��Y��	+�Sg�I�$�_g�=nA�s��ߞh����8]�xy��f��u�^p��ݙ=X0$�C[r��1��y4�t-��{j��:Ԗ�Ƌ)A�<��&Bͳ��~`�b̀���e��&�b�o���?ۆg֯����R�QT��E~3�k ���=[6#9Y�$W���f�D�k^�(�0m�)�]64���A?|{�3Z�M݆>&�;i���9u�ȿ�X"lc��2��N2	��Er�x<� ��p%�;�&�B)���+�DG�LU��a�K�Z=�*��Y�S�
���j|r�7�Q9_
lMu���'�|�ղ���U<p+���ߞ��k�pZL�O�2Ug��}�GE_[zW\���&^�V��)�u�
�Q��6$#�U/ű�Ҝ�q���:�=A�* �;�5B���c���8�\�2�O}2�\��hb�3�,9"��f6[��X6W��4�-ͪ�u1>������G�?Ggfe��+�{�^Wx  ~�qu_t4���ÂRm	�x���7�� ����ƮrӢX�|_x&c�������{�wh�~�Y}eJ��ÛR�nGP?�,������ϩrm3C^o�֖���h��/"���� E��z+JM���<y�O�"����
02}���B+M�4	A&����1��H�0�7ye8E�e� U��������H{p�����Z!���lb�2ɒ�jwo�P����a���ÏjCO�fI�3�O%�c�x,%�����V�Nh������1�	�
[d%}���.���Z��b���!�lQ��YkU���ِ�T�`��(���-�J�T�v���a��ɴ�ߠ(�_=4w��6��"j�p�3���Q����C�l���F��?��>;`.�����f�x���E<��Q�6Ӆ��C2/QT���K��.7A��ى�{K�=)*�}�]��	[���z~'A3����+�@�Ĭ���d�_ [��Z�$}��K�:U�qW�x�!�i�x�p~����g��dG�U޽���<���G��꭪:,���]��
��[�����%�)o�،b_M�~�?�
�����H^��2)��Y?��6AE�։H�)�B�pה4c� .�X�9�@Y��