XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���F�a:F\����H���H�5!$f���݊j�t�����/^���K��≑K@y??������(I���{Ѥpq�<>v?���2s�+{+�Xv��?�G8*A��ɫ�t�dS�|�\�d�<��3l���_��q��?r��%- Ah	�z�+寜L���iҴ��Cs�S��}�~�B�Pރ�ݙ�;۠Ho~V��F"�)"au���n�E��&G�gP���Ŕ��,��Y�wH�����Z��D?��>JzQ���N��"ot�:&N�Ӈ���kn%�ڨb6�x�x���apw[��N��sq�ʜ�n=��<�`���r/G㬻��CF� U���V[HΞ3��,�T=I5~��gL�3�������:��; ԃ���+�e��0��1��r��T���'�:�V��x�р+N�\
���a(���WBX���o��9�VW��=b|4�~�ϥ�)3�Su��kX��}(�1�8"����L햝S�����}̷=����Nf&����7}����$rq�[�n<�ׄO��[�,��C���KASo���t�1��a���(e�Ci�ScL���Ґ�L��7js�f���%yn�+�43�]u��"ж��ؐ/L�Æm�����(m�)v1�,Ή
��L�����$��.��)y����X�1	'��A@/�Cոj�(g���|L�/b��I\�+t����gl����Y��y�ά�֪8�'7����O��ڽ�;Y��2O��XlxVHYEB    4052    10f0 �l�&
Ś1���k���v���*gڏ��<��0y��Kj�_3���۾�|�H)5����;#XQ�s�#��=�Ɠj���kز��΂�]\E_H�S�)������H�<��d&�F{fO������Ľ��<zھ@d��8�am)h~��@�!�S{�\�8�:��Y�|��>.�Y��T|C�4j�'�pl��������u��q����,��F�`�aF�o�!\\0�,e�?�v�*|�Z�_�/M���=��q{����QM洇�^�������Q��p-�����ě������W]v>T�͆ߛ���^��o��D�^�>����ѕ#���)(k��g�����֧c���3� z1*�ywL��cF�[�Xd�A|C��!l��؝����J�ؼ��X����|�����v��iƨ���Ř'm(�m����� /I���ݺQWJ���xHn�z�0��{$SYm��%/��{��?k�?TP���0'�G�
��J����!�12���E��Ov������E��=�ӡݞjykx�C�n���"z�}#�>J��-��;G�`[�=�joe��}؃(O��mE��TD\��L�{���>���:0�)�9�7����_�e$B�׎��j����/�dF�Oؤ���b���Y����rA��u0E�����i��#l�JC�ٰ�T� D������}	ꖸ��#������)�H����@�3x�Ah29u�Y��<�<�	�#-���� Ҩ6�h����?l�����E*&�M�؎���T�g$������eż��tg��ࠀjՅ]JM�i3!c�g�p�K�U���u�}�v����g�JN�<�t	s�hi����}�P�6X�]�C�JB*����Qv��������2�e�F�~�;l�"?lP���9D�G)~���?��WE�i���zVH����F��-�'���ݷ��x�Li�f��!���T9מ-�p?�R�ie017��}�o},���*��B?����:�ZfM�ю<�lֻg�^����d� ��0`s<�]iL��j�jRWJO�qˁ�Ys��f��*S��n��@-ڃDx
�7>�sj6����5�>oJ�E�μ��B%-�3q;��"31�}Y��^v\3������A��c���J�X��T��~����7R@(5g�F�[�lz9�.�A����Dv��ֈ�0��D�^)�����B�y�i���˞�:B�Q�G*gʋ#i��kv|^ AO���w�_���q�c������rZI�Ws�iK Y���kذ���ř���R6�rQ3�l���ʷ1���� ̮��� yag_vb&a1�a��K'ƕ
E������)Y��
r�j5��T�"�;�bAV�\&��.UeWz�Z<�ܩ��]sC��÷�)u8�'\���[D	��V���r�g�)��b��t�ߢ�9'��OO.^:�>�������Ɉj�(S���+��A#x�X)��kF"�X��g�V%�{��R�v���x�!�V���Qm��ׯ���+��k6[���བྷ��Q��ox�fhh	@��.\��Y��C��	�-/��������\ƫ�t����Z5���̤��i' k����)�WG�4;)�����,1���r����Ir%��z��B�TM�!��W���$���@��D�!(ӮAA�{��a�u�gpbI͡� r����/6:W^�W�-u��T�hsD8�+;�T����6��(��`�+����S����+)$���q�k�!Q㢯X����sO-�_M�FN{���mP�"���ۙׯ!]��o���H�$�H�l尩6cܺ���L�ŵDή��<;V�v,�k�4��z�:���zT���./��J��\��o^a�&�����b�j[�=wIĀ �!b�ž�����2Ar����ŠVx�ã+h�M�WU��u�L�u�s�u�V��F��sv9R�n鎢����5�=Z%$M�\{�|�}�mD�s��E���g��z������3�T-zJ.?���;%��L��Fdd�lC��b�������]��5��l���&e.�`��Ν�����I�;%�0�0f����3��w�!^�U�h�>�q�ֱ��)錁���`��Ign}L�g��������%~�a��-���m,ز�9~����
��L8��x�*{>��'�6�9�10q%^/2����ܖ��a�)�� �?���W<F�Y��m��v�XLK��V>T�:r3�P"��
�N$)��g����# _&�cYH۹�84j���M���N���;��*X��_�h�߅S@�h��~8C�4�r��&ms�� W���MhZcS=��r��p$�e�Z��H��i�k�(T�I*ȧ>n��J���0�lI!�;�$����*�H�+��AU��֙��B`W���#�I��^���f�	,'Rv�Oqr*^hWV=!���G�BG^s�Lt#��f�m2 Mt�r���Þڃg+���N��}�U۟��y�QUj~��Qވ�="�2�KK_d��`�gm���VYU�M�1��Zq��-}�:*��*���Ys�>e4��>ߌv@���v�׫��M����~p'�2�����2e��=G��x�ϞP�rp+�����j��cZ�R!�Y9[^�ڑWj�����;�1�H�r��6���@3��.݇t�&���Wq;B�w�:����yf�c���,$RȃM�R>A��q܈[I�[�a8��~�T5C���kذ�7�9S��J���Cl�{��r<�^*^�^��e�vK�Q���Α�T�!�����=�Vb�?�-��`���ayef�v�=�Q-A��,�����F\I	bI�NNЬ��n[�-���J_T�g(D:Ӽ�O׎$��	૰4G:4��-�O���JBg+z���ZР缺OV;������{���ލ���ub�qjH�@��z�i{�{�6���a���i)���Z� �8��)�:F��,���(��ڣʖ*�ԃV��[ML�nI9�Ҁ���p��@�,sp!n%i����i;>�I*^�Ͱ�%��lX�g'P9��W�(���n�k6�`�cE���C����a����^$'9
� ��[����l�-�%u�9<.�ˁ����~���/Q8Q0��x#ŹT�@|˖_rP�vAD}-G���4�*���2 �Ϫ�\Ȏf�"O4EE��-�����{�_U)��	�am����3X�T9�(/M��ρ\}&5l����&���w�Jh��-�����.�Y�$�3\�1E5A��U������dMc�,rt<�Mۇ��
��XEk���|h`���|O��m}8��/�=�o~*�kݽ��w,w#���͇���۽�sߒ�N��ei]�nnފ����qez��q���3%���~�m��.���H5���N4=�W�#"x�ġ�fq��?��[���E��n�C��:�_X�~��c�>r@��[�v��|��D.1ܽ�w��
�E��Y�='9�[2��'��)�������}@�W��#��2���ǅ���`�H��.|��6	N�I�V,n�W#�@�b�y�S���`�`$:$���+���J#Yɲ����{P�2:r�"І��6��+�e:vEg�!i���~N!;ۈ�hi9�@�x�Q�������F���P��A�*N�1��0Z���Q�V�ɚ�.Tk����oa�FB����"�g�����ۣhG�!{���u�c O�#�&&*�}�Qd2��$�+F��X�6[��g>^"�#L;�Fm�a�	����}z�5���̂��[����Kq�cȗ�F�ȋ��̾�}�=q�����ޖ[�ɵ�~�
�Tgs#����dӊE\K����O�+�(�ɂJ�2�v_���=T�����J4[׆�e�a�l.[�H^k���p%�x�5���i|�efxN�� m'ς���2���_��@���E�b��'Q�*�{!�������v�]ο�N4],��D��B/��aV�������z��e�?M�k�<��">��>���եR�:O��Ԃ�{>$'�e�㿶��?|��:Ftm2�V����'+�b�9}[��n����+�_��`` ��F�L���9�u0?���x��F��r��2l_�G�A�r��"�
�N(��&!������+��1�Nk�̱���!���Е�H��Y�I�G-ʅ�v���Ǽ�A[�>��L��}�G��~X�t<=����ȎMI&6XE=E�$���<vL