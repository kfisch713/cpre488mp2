XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����.6]l��� e�ɵc��d��I(�RZ�O�$1A�EXݐ�g%����o9��L��@��UIv+<�{,��xs��l!}��*��f��	��Wtxd�S�4�-zMg�ćʔ�P�CM���KL�����c��fE��
�|���{��)5F%}�7�^-��pGw]��5�)H���g+�>�G���^��=�_��U��e�Q��k�a&]u�pQ�
����Pb����n�N��Y�m���!#�ո�92]��� ��N�g*(���b�y�H��S	��8GZ��}���Z�I�~]�Xe��DD�������׫\� h���6��ke�^�y?ӹ05`yBa$���2AӨX��؇ԩb�_1��1 �J�K���,p��kD�P����;
��X�@|pe�FF���q����r��u B8N�ǌz�ݲ��K}Z�)<�	��+(�5ȗc[3������#���lN�dMbT���߇��آZ$�=hCe�K������/� ���P	�%q��0H���pL�P�uTٸ�MYc��D����a�@��+3=!eՏ����@��� ֑N����>y��=�Ԓ��m��K;��Q�@�9vH�O�ovs�+sa�$��O���@D�k��Zk3�hP��)��
}�"j��;���nP!�X�P���!)\w�cX�1����,�Q�΀�(�z�r*
b��A~��QD'|�6dkul�	I�� ��f:��OJ�@����f���@��C���6�$vAXlxVHYEB    17b2     880wr����Ka�"�������6�뚌�p�'l�ehq�=
�������r{D��~��Z+8�݈%���?����i�ԇ? �^&�?s;6����q �2)T	ɚ��h8�V=���ɺq^�)���	�'o���[X�>N�p�b 6�1k8v�*״e�W_z�D"�dĽh����}Ⅾ��W��r,����?$
��`��3D��|��{G�HR�M�*�<��a$?��"q_K��?na���J�w8�Jm\yb<8L�ʌ��� �ОUJ�/�0[R=5?x�,�-D����C��=S�����S  o���7^�v�A�ܼb �������vO��t�W�:�~��^�T�Ah�us�r/ ��o�q~����֗4�;t5DB�;��T�c�H;������_�=���a��~���\���㖄 OicB��+g��`j�)�E?^� GU�,e��}`�e����'�贁8��l3���T{{�+��	Q� �4��� ��`z��N,�1@�ɎF�j ��K�7�%�mA�j���mZ���?Y��i��t?�J)	�%�]p�����}�8w�I�l��E�^�8�Ϲ�%��?�l���|�<n�}宏������_� a�O�׵qdY�>P��;����#wK�Q�2���Ϗ��9���,�1^LG�^����)C�K���`��F�h`f�	�q���Yy��*��8B��V�|m��H2K|J�_���)��=H��9�j�~�	�O�Ճ����ĳ���m1A|�k�I�qHVI����� 6�[.�J�)����d}��÷��äV֘����[�����^޺[�0�!>2��l�_h�	Zp}��Φm>k�f#�xZ��5*R����yVHo������+U6��x�#@�6Q�{	�c�Ϫ���/c,�������y3_Txjf5U�	%�E_h`��:>F`^❴��9����[?V�

��@SDbZd1ӈ1�Y� ��r0�T���W'+t:"��LL�|��<퐝��b�FIy�x���G����A�Q�.�� �wʽ�g(���2�N��Eӛ�cB1k�q�;|Wȭ{�����uϗ�T7P�gaXۄ�br�10�X�,X�WY��Oz��#+]:JNi�jIG�u�M���!�v�b�o J��A�2�R�p+֧�q��6��`Y��,@�{�V 6�3�R(M���(Hq� Y��C�2�=+j�������>j�y摥)�h\����	�����h�������6u��x2G������������D�U,Eƨ?"lQ��Y�pE�	+�Fw��*�����j��quQh���F��O����I5&�܄=&�46�`59R	��K= ۄ����YBl�H�A��f��F���G�׵��s�0O�	%C���W��V2�m�Nؿ��*�'��	e�na��z��Jj5ݽ��D�!~�f�π)ǫ'�9��A_(ji���T��W��@���
�D��=�/��0��E=N�M7��.&m��������zk�It&:���Ϝ��cNqz����_����)7��v�Hu�`�a�O����j��RвT��}��tܱ�c�[�Q��_��ި|��ߌ����bUVQ	���U_B�e���n�Z'nd���<������B!���\~eϨ����2�ZGG�V���W����?�LД1�PK!CY��c�4"��ؕ��m!k�[��d7����D6����̱w�K��N�l���o��gK�n��޶��O��]v��%�U��_x���c���q���ɃkQ�1!��X�T¡I1=H�� -o��?j�����8sH����P��E77JOݥhLN0������#��k��q�x��:����Dƍ.��4�Ͽ�%J5�<F@@��̆>���f�Z�<5e^�,�T�e9~����!���%��� ���a_S2��7�,�׋�J��E���.��ŝ����N�N
��Rj���5ht�&A��KCYsJ���@���X2k`#�l��P���q,5(Yxl7/"���R�\�A�E�����>w��$�MN\�����/�.�;]��>�ڍ�xiL��b���{5G��� �ju+.�h�ռEį�2��a�[N��9p��3=�