XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[�!���-B��V�>�|�
�\pM�Zb���GX��F����D]I;rH~>Mʶ����O)��o�S��7ˀ�$β������xV�b���F��%�����#fE�N�-�2���Q{�64�8.#D���$�C�ЯKd�WC�t�#-�b�ޛ�&BK�+Xtğ��A����⢩m�Fܶ�@Jh��h,���=��x��Ym��Cw�J�&:ￜ5�Y^�&|367Y�7�"�	@�]zq�_�i��0��d�z����`���{L]e�V�)^�55�c��o2�ו<�
��V ��q;%�*pyY�{~1o����0�`s�v���5�<&]`Wyն8,�O�;�fP�1T���Qx2�Ǳ����@;��8�9�ǥ�9��f�!rH�. �b|�V���;8��ԑ�`jH#�&<N�j�;,�\�շ)��2�zJS�R0%�h��� 
��W�+������;��`�Un��d���>��o@��t��2�������������r胲0��R&�|.�f�F��������	u��O�a"@��n<�Z[�L�<�
䗧�M4�vh�����5$�[�hB[~�����'�Y�~:��2�5
�۠e���UZm�1�;�ΐߒ��[�7�[x��x����6ռ���gG2VY��`X{qe�2�ȰF����b>[B�"��Q����2@�����S����~�^D׬�SF�o����#��F�8p��-_8i:]i4M5�3�濒e/cI��hP=�XlxVHYEB    5e2b    1530�<�u�Ғ��ŏ�E6u�,����μ�9u�l#�*9����/�p�k^B��u��=�j	�Mօ[T�Uf�D�s���d�]�Ǿ�כ��5�F⤴S kG0��a�����W���Õ2/�ʢ�������DM�j&օ�|�T�q	���毉���߷^��UWK�O-L!�!��I����n��R��]��>�S���p�]�.G]k��|���.[9"�T:v�QxO�J������0r�M��r�f@�	3(�jdc��#[�y˺�dqkb��D�I��\|'ج ��o�kige�1+qE�{�n;]�3x�^�����s����!�<�↋�+{"I�$U?@���6��n�|�_�48+SI����z�>��r|
��[+�x���* �
u��,�m�%{믪�J�8SIj�;W@�O��?w�%�T�:�1��d�1�7B�^�NbJ��2��9j�~S�DV��$�s�AHc�պr��*f�F�ͭ�h��o����K�A:�I�5;6Z�ot����Y*D �6>�&:�`@�7@�Xv�5�RxM�I���Q%b����7�?]?��L?!��I?��7�c]D��ɍ撘��l:�z�¼+h��dώh�?iV*�r!�'�eK�Sӫ`�	�e 낆e"��t|a�A�MXq��Q�w�Ŋ�-���5��o>�j�x�</���7.������ e�X�sq��<�M�F�ۨ]9G�/�?�����d����M�.p6���}�u�S��s����z�"22�֌�������G��K�_�4U^ �KL9�3�m�uy�|[7m>�H�9�'gu]����9�R��[�"Nӆ�Q"�0D�ھ��U�Cu����f�yR��'u�20����<eQ$-f���׌+[�[z9@�J��>g�!8f/z�q�g���J�U
����I�*�b�J5
���K2�n��5>��ǽ�*�����Y�h�R���Ѿ |9V������M�/�b-X%��\eR��+��������|�Z��'g��)�j�y�"�a���-P�	437�z�&��
��
��6�Q�٪�fuHc��[m�'�v���3��o�P��r�;I�ȩ8�� �M�?�`1ֺ1}E���%o�U�HH�L�j��-�����qŢO:n��-U6������� ˫�A��"N�1:�M�H�m����YTp��lK���wWrt�W4��5%%4���~�($�.��{۾��P*����~�l���2���z��Q���������Y����u��6��jծ��������1�{3rP��YAĚ�_�X�3����; {mA�JIy�j��Ef�[4e��ή�RFrE%��D��Y"��i��&�R�tRU5O,�gz�X�w��{D��Y�;���Q���V�y�d�U=U:_jƣ�'��,�z�w����#�Y�4T@��Рu��2B�"�HM>1;���2�����~�Y!j�E0�f>����L�ע{��!�s4�Zdլς�j�����1����8�:���@ԭ��������Y�6���(͟������2J�?x��d�c'?d~�r�_������,�) U����p+>�«.l�����U�Hh��}gN�kOY�� �s����.�<����B��R)���߁Hf�r�	�w��[�l��wrO�%�1K��gW놅�k.y� C�Wś���ѧ><K��8��\U@�j�"C�A�;�E�$���f��8�0�%�=����񃐙�����t��I<�SY偘�e�RS�m]x�O����=�}Â�QԳFh�X�ejG@4GPF�HPϩ��(�!��iD�e�wL*�Ǩ,L���v(Z�aA���:`JW�� ��_�����4֡�����Z�ӫ�+gA�"FN��R��8�0HC6����T��t��No`���v�ϩ�D�
�ۻ��taZZ�D��=���t)P����e��}JF���?���\�A�|+?נ����]z��̬1��z[v�H1��}��>!��o#��r�Oy��[(�I���Y4=�;b o��Y�� ���,%N3:�D5�o�0��)��k@~��:䵂�84��IYgz6��tݻ�(�nb�Re"h�
B@\`����}���j`Q�[
��-�llˌ`�̊Q�\�b�u���=Ƽ�?8?;(5�&�$�R�����7�;�;���s����=��MMF���wv�m��X�
�`n�z*(Q���l\���r��<r�X��u��#S��u��]<���j����l�3$�*�/7O�E�����2lz$�2���p&����00g;�v>M��Ed�\еẊ�^�~�V�)5R���4D��7DC�+]N*x����9 *��b�k�"�w��j�И -��9�^�7yO{����FWb@�q޹73���p�3<�*�XA�WX>����/���F��Q�6h!x嬖\J��,�OM9����CE�WL����)�p��S{/IY*�r�[-���C�*����?��a��$�(��O���p7o�H!:��G`�y ��\��(->����H��ZHOP��Ky`���w��t0�B���)Í��X��x[9�G�+� �q�@b+�w:+t[ZC2���Gp��k@�1�O��/E�m�=#aR��ϱ4��17��ڿ6C*�~���w�߭Q�X+H9Z�}��Z��ao?�?���j0lqa���~E,c��F�}�~D�
�I��D#[����3j�w�E@�m�\�(����\rĨ�u�����Ev�4���[����w���*���9���U���S�2�ZZ���y]��X��<U�>e����B���y�{�&�J{�K�W��G�ѪI7g���meUP��P��9M����y*�����?���!��S���9� ���sV��NU�gu�o��PL?M�dX�vK��n,q�B�1��CHN�&g�� �W��2K�Ƕ9�)�%_�R/���
r��W
=GM�"p����%z���n�(e�_�{�]X�
�=�QR�H�%oX֞���H�H�J#�VK4���EOP�M���z��X���~W9|�*�,��A��T�Q��k��u
�W�)� ��ަ��a-�>M��|���l&Y.c�6OO(J��4�"�6�ލ� Њ:�
%�ו����B��*�]S0����7kܗ�2ZT�-�BqZKd
�P�/�&�.�lX'��Mr����
��H��Ȕ$K�ʡ`vmkށ�f���L1�$����P�ԯ<���^��8)�<�Dc�|m1�"�Y�E*�WFk�'�ԘiTo�=��G�B��_�R�a��A�\<�6G�z�
o4��,Ō�����y�LT�?��.i�ˉf܄�x��*�G���,��7���6���C��i�*�tNm��(ґ+��[ڕ,˸,�h�XY6�00��uа�W���7|..G�+(�]�g��Jmv��Z]���<�����Ld8�X�=�TC�+��L+���xQbI��p(����5`}�0��Yg`V5t}�m�=��= ��x�OUt�(�Q֮�A+y�G�J�����o�	S�A�4�?�S��M`RZ0�ة2�JE���{��^HY'����[�2Æ��M2��|B��7)�/}�w�JE$�9kfTD�z4q�l���+M�-��.��t.�5�<d	k|�{E�;\�s��y�"�GI벾`�r���9D�h��ϣ��9�� �6q��H#\AV�]lz7�	K[�W`�ܧy��e��x7����Oڊ-�+9�����	߈ݏ6���G<b=W6H5K���E��5b�e�����<]�۝:��>� �Ȅ����?�\	ݑ���/�����B<�= ˿e��UPO����j��7EÖ���f*\����#�O�(I>gD̫���Q'`���P�$L��(��]'�����02���~��������<��R��ϭ��1i�b��l�x�9��Xk�/d\�0|�f''��<����q��?�5�0�'EB�y��f	�PoVaԣ1a{	9���Ap��J0��3�Y�Ƙ2E��b`z��a0~M�3����^�GLCF���W���DϬ<�C|;�Y�=���l�!�<��������6Z��߫R�x�#�� �x���gc��Ϝ�!Mű�8�a����u��  +�r���j���7bD�+�͘�+��c�@�`�`�'���n��'��x�#��_�#�]j�?|�����W}�y�z��͈���>
����⇏�9C)���R��j�����BYY�������; W����%�A�O����*g��1��I^��N�+����ֽE�(,�g�!�3���5�`�N�~�M�~��{�o�K]x�v�Y(�,qcnv{�ɒ�drY\!�AO��r����>+�j_ pw�q�o����K�ȅ!qk��h=�a)���j<��,����#�{���0�8Q5G��Sq�����ڵ�Ck'p�ut�~��<'$���g��uj��p�=���tZI��Q3~����!�3'��Aw\�"b#b�c�������� �E�'ԄO Vaw"�ly��b#�1a�u3�O��Pi�͟gK�<b�N|)�r}TvlZ��%����ߠ1�Q~�I%�DV��V ���qTMJ9������&�_�g'^/<w4yN���ų�0��,��p��F.�f+��:�R;�+�iEȝ����4Yb�;������Qwp��q]��^g{H�A5L���&�HҎ/Dy4-�J�F��ꤼ`>"��W�>��
���-Ð{��%����Xg!c*�>�E6A�7ni]O��`����޳����m�8Ӣ�b��xͼ!��xה�g<�t ����gB��N2��,� �Wt_�桏z)��ȁng�#�e@zcC��lɛ���|6�
0���B�wS���!# �H
����v�D�����h /��_B��ɸ�����-1"�b�T���St'@�0b�CR�:" ���P٢l_���'���_�}:R�Y�~��������ACe�����+�=����~����!�Q�51s�r�*DȠ���j���#s֗��M���(:ĉ���p�8pM�ޚv3�\�����:6�1�^��i����o�O4�f%ix�kZ"�I��M��}$�|ﮨ�Ad�y���t44�#d�x?��I ��"����л�`V�7Ԣ��@�(JK���Ϲ3`D)W����d9b�nM�3ц����q�=��k�� ���P�� ����f��2�tv��?���k���ԌU$7?q�3�������٧7�)v�`��YQt�ۦn�