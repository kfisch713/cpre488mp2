XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Fpkk齑+M_�W��A�ۖ���u}V�FH8�k??e�Y����¸� O��X[_E�Rk#�ݥ-}����@W�w�Pyfy0����"�R�Ռ� u�2_"���0`���o��!�[��]�|ҟ�z��V���I��Ə�MN�[:��U���V�5�	��Z�T-�z����1�OH4����Z��K�]��Z�C����r���ws�D"|��T�d�gz^?��Z�JF-�ʓ�� 5iu댋�B���Tm&���χR���	�tZrW�<�� ,��^��DW�]1~�h��n'q�T"tG�iD%����]ZVI�8YI�Ľ���c�(���ʆG��,�+�`1$���oz`�v��&7P����xwdd���p�N�8����.�X\�zȤ��N�E� pO�X�A&0�p��� $��ϳ��蠁��;Z?��=���Z�iP����k
��ѐ�hs�w�@�D���?�	��r�� +�W��y��b����Qs*7[��c#�{g[,����/�C�1F�-Yy��Ndu�@?��.�+:�!s9��p�b�H��0#:O�E`rn %�rݩgq.��YmF�f�+���yA��(L��%N��Ȝxh����XBY���� ��W���+�^5�9��H@�X�7;׼HQ{ą��[�Ğ&���t%o'�K���I�F��:nv��'��w �-o3�т�X�@A��h�-2�j��/]�w���
�@p��+T�A"d����[Z>3��e;�\��XlxVHYEB    5d29    1390���ʃPHa�|�^`e�x�\����|�Z��7Z#�c����gn��2��}B�n���$M)��N���fy�� ��V�a��s�`�O��f�4׮�
���Mz|��g'�<Ɗ����6._����s�y��J�5�s��h�Ci��!6 짦1Q:�1�s?����pūk���$��: ]�!�-��@�;l�|?FI"|�bu��q��-D�Hv-o�0�q�ѩ������:/{���6�Y>��wB���'4M���P��|m`�XF�p|1�Ŭ1�R�8k�����w�Ԗ���8YF�/`>`I�E��x������$�+�߭�f���Q ;
�Qb� W�� �#�N�O�2����� ��R�T��KlC��o�<�N�jӲ�Z�^'Y�����<Ԗ�nZ��vV�i1C�佃���0E�jl����3�i�����S0�Ɉ����[�x�%�;\�1���0:��T`��� ��L��0P�x.8�i�)k����츪 �0�����@�]��M��ze)P���qߩ����R��#]V��B2*[�M���:�*o60[���C��lA���tb`�-r��q�M�l�D7�`�HA6��::B�֕u��[O�Yl�(�(%kM��p�5��1���^2YV��������o$D��ܨm�ݡK��˂�m�_�o�_^�Kk�#F���٬����h��K��|�!�"V|c:wi�h��;4^�i���>0[):��D�1�)�hTC��Gu�Ґ��)+��%}��7��������x���J�h��;��7>]��]�����w��n�12���f	�h���t�ޟ;Є>��2ʔT~��M���Z:{ụ̈̌�Z�8�(��Sx�-H���f���;f�+�ia/�f�X����fH��k�i�!�4c6_dԅ�F�6�fE�>)VT���T]��,�#���
�����6�0�{7�~;-~:LɄ��‑k'�a�v�����X�5&��w�{A9ܡ�O��l������l�nNr�l�c� �!���8�r�	>�3yS�J�9�_�Z[
�EɍWv5�[���]@i���ؙ?����6('f�F �/�+�H;��`\�Կ����暪*�/��=,����IR򫊩�����o7�2��~m9�k��0����2!<����z�����Ag�|ơ�>nOMފ�^�3���S��Tre��z�k�D�GY|����&NK���`hfj56��0��zW:9�]�61/K�p�. ����'cc��J9�.Γ����m ����(���Gr����0ߴ^g��ϐ�X��p�L�/�o��)ڤO��ih��w�aTjg�_>���+�#H��Z��z��M�
-]��sd��>� ���SХaߛ�6���v�]��D�3��9Ԋ���߬d3N�1`� ��Ú�^-Z�5�H<C�|s>Og�8e���~�0�d�Gm\ =���h��u��jN��吂ݕ���T��#�r�����n�9b|+U/�]���$�ƫ����Lc��ߟ���G���aq��Ȍ���7�?&�".`�݄�B��>�"��I���]n.�N�/w�X:��H�$�E-2����R[�!��t4�
������[؀��\�*��9����������Uq��\+*?�$��������e߆������&KqK�(	��*H]�n����Í5�6M��R�������T��h�̊��&[&d��`���3���`o�?��݆���oPO�Č��2����
�Ԧh/a�w��Ϡ�o�O�qf���61Go�a�0E�4<��QϢo	��rh�H���B*]������I�rX�Pl��dnn�~�z��{�CW�[qu��_�甥z�J&�G��(�:�bXG��w�t�n!639��mcȺ"0ޣ�T�ՠ�7UΏCx�����ބ�0J����Հ�����~�f��@��0`���%��[%������V[i3A�ZϬ�8N#Va^��A�8��(R���\n���w��ヿȿ��ASJ��j���"Q��o�rgSk?�d��u�7vՉ��} ���w�����P���Hc��|&>�:�@�w��B������/�t����{$3��hL�0�vt����;����f���p��Q�o����[�mó��"ד�I�,89ha�2�J�T�"b$j�0��)��*�xp��Ny�K�H�a�XSc���?L%x� @y�/�/z>gu��DQ�zRȀ@5��΋A /�Ǐ�H���dV���	즰�p����S
��7�Là��؉/sYLUt����V,t�{tfw�BΔ�_̘����h>��Tg�����;#��AyO�>z�)W(}�n;_���A�N�B/x;{
T7ΨY?���C7�[��P�,�><�7�y﷬�ا+o�wžXvG��v�B��¬Q'����ϕ`I����܄|�	\����tU��e�Y���������Ħ@��A��g[�yvi`p4ב�&�n�r贿\����`�?�*���g��o<���tk����n��r'F���	b�S�!�BZ^[<,4MF5����$]�29!��ב�J�3m�S��[p���8��!_ ���dw��L��νalM�*߫N��,���:�X�~�C�l�Y"=v��k�{x z{֫�����8`�%q=������,o�}�(/ۧ.��?��+X�#�hv��a�İ���� nXCZ���2�(��5�۹�����*�I5OJjHiO佋?pݴ)���:��~_Bܘ�?�ó.<���x����򝴯(�w�N����i�y'S��6�]������#eW�����n�����h~s��n�!��m\׃���&���I�i��%���ޕ)W�ך�������~���u����gV��8)��ɽ�l�r[5� �Xg�x�7.�):��8V�����`i.�P�2>毛&@�V5%������\�E�c�'潦��n�x�^ 3)�����Ĳ繍�ѱըbg2v%�3��@Z�M�j���[J��>���6�a��4�|]Ĩd���#�QY/��;�c��J�8v����JP�.^90Q�� ���`P�:�^���S(��`%:v�BP6�i\�'�N�/s���Кk	I�C6�k��|�ȯ�U;\_��H�ll�
���Ñ�k���Ҧ��Y�Uz����Í�V����p������ȍ�*P[��Y�q� �ѡ��@��L�Z�.���MP�e�� }�v�IT`��e�j�_�턞��<�xP���KSA���fԱw4F���S%����T4�]�Κ�e�R�J����vS�`���j�_�z��h��]�}V��k!:�Yl��e@��������ѳ0UQ��1��$x�*�K�$��F�|�Dl�	=��ꬢ��A���A�e��(�dN̸o�q&/W3��D�/A�?0^N��\r�f��L_��#�.�*�͢��O�0��C'�����3g�Aoc�iEٺ��R��`FI�5�|�k���p<�h�j������/k��+��(��6��.)�SK�C����1��
�	l����qy�긒 7vxC�8$Z��:���2�#���q�f˒�U�K&q�0e�	��P�r�y��>���y�+
����w�  �9�1��bfkt���	�֋��Z��YJ�uԩTY7��rn��d,,��)�<.E��{����c��fC2˛��z�1����S���T>M.Z�79��}�m���S�uw�3��t6;1|�I�" ����.x��vA|bQ�� @�x���{)�G�&�}�%
���Ȉ�(�=ɥO�'0G���^��� �"���S��"�wћS��4/�7����`�M��Y$�?���]S�XǄ*SV�%KM�sE�C @�l]U��w6�IYu;q��醕�Õ��=n��H/A
[��HF(�V%�FDR*����3e:31���Mz�� %�%����C]����X���-x- �I�/��B�i���]j}Ĉf���^]��f����5�	A�S��:.�ˉB�� O;��s�4�Z��k	Ci��4V�<ě��p�����K��Q�����L�q� �1�,�%��k�����Ĺ+/#�0��=K`�T��)����/����Z8�� ���i��u\���[K�9���XB��~�twmb�Z�a���Cd6���GD�?g�.�0>I3�Q-�}�#�����,5�!�O���V��}� 7b޸�$�d�r�
lw�d?�Ȭ�4�2��Ƹ?O񿼸��>v8��7k���?��9E��L���| ����m{b�5.������eݰ�;Z���҉qƉy��`n��IxԘ��:�������p�-�n1����겚"�è��ݤ�{j�|P��G�l�>��
V5t (Q����߰@闺�w���&y�=�A88~�!*�Ps��e��_ �]cq�N�H��.�;�s���KH�p�NF��5�|�+[�x����=�]#X���90*^���� ��2n��',�� F->^�l�˹�}P��ˤl�	�k�#f�|
 ��$�5�4.�W��x����@
�r=��@�&�v��)N4?��Y�P�J�RւGZ]��=�|��аR����4�����W�e���捄�Ł�l��mjWoz짯ƅ�����B�`���t�h�8q�l4�t�j۶�[��C�q:���Y�@W:չ��kϐ=?9����kw���u��b&=W˜��8�z�v+Ɍ��R�߱õ+/����V�!�]�X�D�|��(YK�(Jc�T#���h�o����lG8�9,�_G%���߂���K���b#,�����e�ɲ�O���r����Dq��B�6X��*K�DI~(�I�U�����, ^�MG=�\E