XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@�!`��cm�J�5��$����Y���I	�F*G�y PH`�K�V�_k�Q�q��$L����Ws^h�e,�;��@%ē�S��˹��@P1F��H���}�R�������B���X��m��nW�E�Sq|`:g�m� z[3�_���{.Anw:��Q�بa�'H(��|�������$�g�|�5!ºX[fTWI�ձk�#2����ߏ�l�=g�IWE*�K+���v�{��Z ���J��b�t9F['�4|1y�1���b�y�~ �v)Fo�o�+ƣ9� (Y��64$�}j� uO��0<�-3��R���E�&��d�b�U�R���*O��z�_ȯr5V��@�s;cF�9������	Ghx���ܻ����$2�4�`�y�x~�������.�ˁa���Z>�g��s�v��u�e
9�9�gϗ�E��U�o�^A	�"؍q5h�e��X���N��*��8{���ܩ�Ӧ�vS�c��p�"N��1��r(1��e�->�h���T�Z� �)���к��LǓ�"UM��L��T�A%L2Ɠ���]�#�.u���ǻ�`T ���t/�v]	�.e{B'�х�y�m��z����I��*���.�\-n�<C�T���FRN���|�@ʶ\��-�%L�e�(��t�q��y��mャ�I����tbDx��>(��u�A��<�S(����~_⎈^�Q.!��_g�Ӗ�926w)"��v⠋��XlxVHYEB    5fea    1830=PJ��� $(��]��?`�3s�B����>��4�[s��/.��"ǋ�������������@A�B=j91�0��Ӟ�f�\�V�+j��/9й����䯷�Ty��H1%�n>S\(�s��HfJ��*Z�끕)�8���l��1����.�D.��j� �B��r	�7,��b�{��P�Y;�����~�m�eJcw�����HY9�T&j=Ր���	R�b�RF���d�"���E:�b����Y�@�������U����	n����o��1�o�ެ�삹��������Q�7�Wa}xؖW��!��%?�I%��A�ڎH�nJ�N���tȴ��d��
�)AUWu_��.�忿�e���\:L:Yϗ^�H��U���W���u)�	�%u3b�5/��3i�o�s�(io� �0�Iڳ�
�۠�9����|$�"#,��dYK]��️��raB���b�6ř;Xl����I�mf��:\F��==Do?^ߗ�ˋ�+��ϵ��VL��Q����*�I�Q��Σ���R����Z#���DO^�+rԤd>#�!�b�v�B�:�x�����\��woW��!�-�R��VCè����Č�X�xM���Z�2R�Bq1�E��
��e���VuFگ���֎��ER��0<.{$ݦ8��
,2������2��u���@�_��Q�z����P܇���m��ȴڮ��� 1�.G-�n�������&���&h���Ea.�ނ�ɵ��l�t��/�9��۬ b��4t�+����¦u�!Q��ɸjV���
���v�$��h7��J1E�Ŀh�^+��uT���]���"e�{��0��}�a��yй��X��_�K��|NEU�@��]���y!G*EsO�o�q��ђZ����8�̥f�ro�����`�.{f�xɔ?G��X1��I�Nd��K�x�һ��9pE-l�۷��?��%�àd�x6ɺ+"}Ih���K�Y�ܓW��p��xv��׬������{7����~�{�?���
����c��Jw����rF>ʘU�tLs�hڥ�������X^�qa���9��&�w�E�M}#6J�����#�iSv�浉�.�e�:j(�Q�[�┅�ƽdI�~�=7���w�&�=N�&>@\��1T��/�"@Twg�ķ�U��)�2�ه�d���ZSc~�������.�)U�l� ��|2��ĸ�S�.i%67���=���)��}hN��nG�6��ʨ�5�U{�5&V�&40,��ۄjB|��0Ih��L�a=�lx���^,(��Y��)���~/���2�h��Bͷ��ZN`im����e�x�T�ZP�E��VHc
�/`�pm5�e�)N\S�����f�CG�vG-� '��B�4�I��2{��H�[��/���{:�Fk�,*���zy�9�3��!�[��bAf<�#�{b��}o�{��w��%f����ϧ�]���8�%��� ���!��3�+�А��a��z�P�[֏�� ��3`Җw��\���,�l��ϝz�
;ȼ%��r���u�P�Y�5���V*[9_zy�{���fF�R��[��97��Aߗ�n���[�x�z��-X�|�9�Ğ�r�X\s�� �$����g��-��҉+��ve4�_倱��)_7͵���q���9P��p�=���(��*~�oaG\��N��I��=s���r�|l��)Y<�v��Jn�u�կQw���fR����B���rЏ!��
�`T�}���a�S�F3�������q|L���"k�l��jb2C�'�`eŚ�MkH[.],5��o]	�4�1>�Y�w�+�1�CudC9��K�*�4ӂ�F������Ob_�׭ND��B��Z��hk[�mb�y���B�Ұ�jz�xC�����I��[�	��.����fi�����7�4��dy/�����_�<=���FW����07z �#�/�<�I�jDEs�Xƥ�$��",{5!��T۟�㐢}��)�]��S�"�w� E5�^Y@�<74LN=/Q�8y�z�ľ-���/���Oc�A�~Q�s
�V���i� ��n�unz��"�����d�1<?4��gPn��A��F����X����23PB������ϲk2O_[��gT��U
5ٚ��iTM�����|�Ps�-6�t@���ޜi5�/D�a����Y�@-��T�*�<C�`�	�V��(��LL��6������UU�`5�<K�\��Y{��]l�pg�/ݨ2����I�%��
�����j3�W,OvT0��QZ�%�z�ߒp7_�}�T�TP� �+�i�6g`�K�ֽx�UU��
A��4��+�H�0�B��ðP2*=�dZFT�^sm=u���H�^�uM�
�܍zs�lt�ZS{4�ZYe?�r�H!��;͐_��C����<�	��$`\k�]�'<�f!�����zE���-�G����eg�@%�|!	=~]�E~��@���ΰ�c^U�v1e��g~��Ċ6eZ�8V9^Wr:�~Co���z��z4���V3��O�`{{��^�&�k�r�Y'D�Dp��\7�2�a�\F,L��A�h%a�\��y�d$��다>@�����␠g�͋ݸO8�L���}�Vᑘ���7���[t�ݶJ����48Т	=�薂�j�;pa�ǜU�_�n:
���k��?��B����#�hr!g�e;���$�����m�LمZ�YrBܯ+]aa�iސ�Z��o�Y1>A����q��~��b��C� ���
x ,������O��`�΢�v�ׄa� �L䮵���ᔋy�?f	��]BLB����wh�,<�Ty���H��Z�iQND�i|�D��ff[g=��X8��������ݒ�!�}����r!�Q��"��Sf4?�ȜOI��+�fX&o3�� ��j�cR#�w�H�f(����,�Bv)��|�(��x���.#՚���Q��/t���&\+v���'y'�m�h�4Zߪ����&�bM���Xi���C9�yR&���)���%� �$�Θr�(���`�+9�*�,�i��`.����F�^���U��Lh���+Xź�\^,F���i@Z�Ab���m �@a�U:.s!Z/'��>6m�\8Ǣ���k�Zkѐ��۟�!�K�������g
�pRS�T����0~�(6�p�K���Q��ԧAn����9� &���U��f81
�Q1_������m$dx��w�H��9�Y~���"�A��-�s4̺�e��:u�]5n3ݑ�c�&2AY�$��F��E&Vۆ�O5�7��g��2��z�r��&���|$-��&8��/)̴<�T ���ba,9`�Зix R�N=ɾZ� !�q|ڋ�/�����ڨjAGZ��6�.�NY�����1��[���F�-&�pk���S��<2J��hw�����U�f�6[?�� :���F�����xpV
6"��LN��+mF���E�Z�W�7+����2!��KT����D-�X6�G�!�s�u��H\	���tG߂���ig�P�6���m{໒z�:���d4����WC�2�ֳ�e=�� ��B&/(��zhS��-0`�	�U��F?|_��	,/����,l����}?�)��%OE�S�S �ê�,'O�����a6��WY�o��&M�2�l�
���8��q4�D�4�}�4.D��y�֥�(�b�%��ou�23qU�vi!l����6�! �$M%VL������!�5!\��l?y�|!\~c�HI��p�&T��X��ڗ�\J� -�W��A�r�v�r\q�:�DT���%�����%�R$��	������G�������@�V�WZ�����d� �r��@+�@��2>�BJ��G�'	>�c�(�ihbz��N͎iB�Z"g���Gx��u<yk�8#�7��e0n��v�7�����cR['�����f/�1�I�&i[���ԥ8�c�q�v�����tw2^�Ze�S�U_4��(o{y�����LxU`�ʸ�#�i��]7��;�_>	�D�"��� �����o�Y�-����t����k��ξW��IP�㠤y/|��:ݭc�1�_{�/�=Y\�Gs�-�[��u�ʝ)$T�U[l�p��|���Ĕ$ zI�a �����oa��%ߌ���iq�ߘ���)|�^ʴ��lY�݁��h�]þ:@�{��?4��
�#��BId��ߜ�C��Y�?�ttz�2�ڔ~�l9Feϙ�#3K7�}�~�(�6S�b��G���X���J@��y��b�z7k>������~S�]M����s9E\k��0��n��;Z���R~����r2T�2gC�d�ֻj�'
�v���Z=�p�cU鳯C�atvl��c u�<�����N��	'ͨO77���,�HP�
���qY�©Td:fX�噴u ,�.Cu-H��;`�N����X�9T(�&�����$I��Ӛ�
�T$�b�8lJ���m��ڑ�XsЊ�
l=,�V��kS3V�:8ݝ��C�l�J��I�^�����d���@/�� 7��N$N7'��5Հ�Fd�u|t7!�#��H�>�1J"�%O�B�m{8�r�6�nK!'`�I�̞l(��I �6�Cj��|t޴ �&NE|ɉ%*V43�0�ѩ��;��e �&,���gqo���/
<��g���n1��nI�Yc���2W������
�K��&��b_8'E��[M�)n/�$�""p�@��9L��+�ZcB���w�5�A���	e�
�a3(o�z�_9��x�ۚ;O���A ���"��[�W���%��$��;��B�{���$�m�sL�	�x���6
�}��L�r{/OC#�
���4�����	{5C!%d>�*K��4I1(y��)�8����\��?��ۨ�'�o�Tu�ӣ�4���`�}�HP�>>GV��x���8 �������=���_&�( ��բ�X�����?{	����He��.(v4��H?��[a�`�k0�5]��X�'���i.,(r�X:WR �d"�.{Iz����K��Й�{�l5@ ;!��ZΊ�>����*W^	����Q��� ��^G���pp����LE�� R����~TL�H���<i������3;���\IH���\,�PU������s����>��'���h\|
"xԕ���Wmx,h]�i�*)�o�|�l��Y�Ɠ��>�L(�M������s6����k�����Бy�����Ú[�7��u�TL� ��VC�+�,2vs����焿
�	^��[�ܰ�{f��3#gU����#�hb=I�Bm>��bO���ؔ��1�yX�P�f���0
'���p� �̒m���v��,;dc�N0��|	jC"D�E}���;��v�P�毟H-�?�ޞu��ˏ�(GbD�@,.z?P'�0�g�Рm��]�����;"� ք���f3y�����I��XhnH�z3�n���2��k
E��7���"qс�Լ�aD���:�!d�a�)"�����Q�y��^_�h��\�MF1�;ⵅ˝�*�/�����պ>��{�P�*�jm��N�&c�D��S�Dc���W!�6�sx�'�A��"+AO?�5��f����rݜnr�4��Ʈ�i/�f�@n�[-�N�W�c�r� wFvi�C+������gP�r���Q��q�Y�����*%t���=W�T�l�T�������k��r�#��dz�'okq�O'�����߹�,-=Y��9Pu��k�hS ��5��V���08���uy�RG�@�?��=7o�	Y/)��'�*���]���1�����C��[8CK.�T¦�����J�*b�v&ђ�PT`×�O�H�[f���I�2:whI�Y��
)=>@4�sq7��ڼ����^xx�cK�
v��o��<�oψ�S0��.G��<��­�ͼ��\&7�4��/Ɉ�}I��Ay VJ�z�ʄ�g�|�<Ϲ� ��W�A�Z8".�6McȲ��� 9�mn�ެ%x�Z�����P*05