XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>*�t3"v���e����%n� ��7͐�d��m�mc����������4�&�@Mif�j�]�z͖��m4Q�8��ܸ�m�O��g�S�t5.A�K��/�*��T��1�4[�e]�Lf|�ZL!r%-7yXr�3 &y�m7?$,�J Czp�L2�/.S?�H3�а���>�E[d����e�y1��4��w���+_�o����f�I�{&��NEb�'.�Omv*$_S�
�T#z]e���%[�l |0��c�5�ù�D �z�	�W�1T6�(��qz�a��b��s��3Ey�DŻS�̪3poj�Q��+z���x��T	�'��Jd�ot"������C�)�L��LA��9�����I�������c	-�<|���Y���� 2����ţу��v��M�{	��d*�s��xDǟ$�[��,�z�8��Fh�m�GD�j���`���zOy��\!ĉ+���m�N�}�Z/Z}#���<� 3ç��H!��s��;�����)&�!a���<�%�<��g�.�)��NY��8j*������Pj�N��OPҩĝbxI��f���q"Ǻ9cئ�Z��L}���I(�(/#'w���}1�x
������Z��)�o4b��Χ�R�݈j�Z��r���ۇ���M�����G���Nތ����7�1�1���K�@bU@+��n5�A��ۛ۸<�hA��s��//�΋�EtTĪ��=�f�So���2�f�Y�1gj(`�@[����a ;>�nXlxVHYEB    1853     810	�K��q�i�� c�}s�]�-�v=`ɮ�R���6���Ů�텵B�
qx��B�/Q*�d	�E�!w�뇘��_�E������W�%��������77~������RctT_F��0c/�:���|t�7����|���C��d����J�Eۀ�$K^{ U�S��Êc\tU�m�BR>u[@�-騡�7M沸�,%��!��
k�Y���/�E(�W����3Q�yUxm�1�`�Y'�9븟�jtD3�M�$ľ�GC����jiU�H��<����-��!H�b#�}��P�{3�|��=�C��� L\r1����՞�ܙ�M���~a�o ^%���j��CI�x�T	m��}x��L;"�ڼFe��aԸ��x��4��Q+ 1W/Q�
�����볽���M�� ��2V���r�AV�)ͻ�U�]�-Sy�����<�H�Y���;=*D2r�VI�$0#����c��i˓{�����?��/@�ղ�c�p�ʈl� 1����Kҩ�q���E�P�+�y0Ң���������=�� ��!��㢓�%K[-�M:޸��_�D�!�W�a�D�Fm����<4r?�Z5o��7���- l���r�,g�)R�@�}�T���50|�ݙ2�6Wy��������I�9�
��Ɵ}h�� ���J�&�%����D���o���a|7MpJDW]��G0_�g���Gγ��Q�����ۡ�* 䈷b����f�z&��i?��0*lP#������9۟5�dƂ�6��N �E�{��X�K�ZZ��fW���3�B�:@���l*��t�}2�w�k�*��U���0��%�+6��Y���%���q3���%͖DT';��Eq�W�(��ޱg
;?] �}&�W�g�h�r�p��{����,'���}�[]��E P��;�h�VV���	��(����o<�`�5�7ss�<��Sq���Ҽ�}K
�*��fpX�k@��+�6�؎r���T�&�*.�S��Ι�S��$����5������Z�$E��t^��:4��4���M�!��)��w��z8�]�(2��/}%�	��h!Lڙ�)&3Ŝ�δ�Ֆ�{�'�iF����>�̖�)�l��«��X��ӈj}���_/1A�'�'�0�g�M��"��+�H%��*;e���D��D.A�Y���z7�h,*'ЬOA/�1�m~X���D�"�4W&m��הn��ͭF��m��tO�HS��V2���ao�]u�} 3#�6�/���`��}g��/T�?�$Tto$BY�8�f>��UYL��h$NKo8V�'�v�1�I�U��b&�&�%������[�MV�":�k�x���:_� rMO��� �Sł��DO�W�H5	�#5�kG�NP�-�����FkB���ِ/�IC�* �C��X��8�6[�O��
�*kl����
�LQ0PQ�
�x���_�Qne�J8̼�=H�L��Vŀ�����0.�ŹA�^�j���!�%�^��bǗ�p��r]�]����7U�`���>S�G��4��6�:�C])�_����ýĄ�|z����������g?����BZ���J��K*g�x��~�9��}����q�A���e��p|���6���J�x|f_.2H�C
|���6{�)>�O�t␕<����*��*1��a�utVA�Q��_<�� ��\jyc/���Å��W$��Bz���_U�y�␨�AQ�6����g�)ĮA��� #>��qG�|[ʍwE�r��m] �0��
mpP��%?h, Z(�P����<6g$Ǡ��Ý��q�a�G��P�w) _�Ų�`.�<�!�ԣc����	�*���/uK��6�̲��D1L����SZ�7��E��z\uM���W׸9�Z`e����"B3����{K6�
8�Q�0}n��L��T��0����[�^��;O����4�;僀(w{�I.y���8��	�EE`���/�H�v�GF~�~ӚO<�>��4�%z�"N����