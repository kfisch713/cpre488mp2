XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��QT�-��8/�즮=B[���dtY��.��+t �P��h<��q&u��l��}�Y��iE	FOn���p��,G�~��51���}dU<������׸$�X�l�"�h��h�oH] ���
�����]��!s�P>�D�%]  ��.ٜpN�1��z.l�W��N	![oL�`\c��)����d�jӮ&�֦�z��_^�&��x] ����l�����e�q��Ðt��NJ��_��R|��\BW�v��_��	j3i�>�)|�H qr��%/�ˇPA�I6n�3��a���,K9�|{[Zj"�����	��;]+H�׾$�n��p��H�x�-�U!�
USEq�C���L0(V4`�8�.x�� �CVl{�`a�4m��N�]V/I�y��5��ؽ{��4�

�LӁ��xi�^��[)̡24V���^x�h}�$מ�!N!����un��U֕̎{^(�$-;X������ �B\ �zOp�΁�j/#i��	f�qB���M^�)
P7����TY�2�(�6�'.x��,���Mk�̜+��J�^�z(��do`y�܅�`�ogJ�3r�ᢻ��l��ۡ���DP���4�9���\�����2c#��9���	�3/��U,�-ݑ���,�����6`��Q�g���>`48y��pT���EZ�m9�s�{̈��nz8M�-�M�B5�j*��Į��:�����o绿`�Q~M���2�>�tF�9�?*XlxVHYEB    1853     810�|^QT#�A����K����/�uX{]�9��1��%"�W���d6x�<!�������-L�K����� R�׎K��UZ�J�6_W�K6���]hf$Id�ߖ+��l��΀�~�2�)��'mh��qn:�n����e�|8V��6M��=LOq偑4o���PF|ت�*+Hޟ;�
�������X��έK�m������A�L��`��QS�&$�r2����b���1?FfMN�����Q�]b�L��3��k$�ɚN����-1��S�,�OW9�d�~�c���xŨr*7�%�����Z����P�2���so�.��X7�|m֨�m�b4.�bT�z�=��b�ݭ����QM���|?��Ŋ���ó(�B ��
VD�8}��f�D���D��SZ�y}��<��K�Į.��Ne4K�nݬ{�[a��8눧=���<�4O��(�����k%���C�n������!����lB�ƘBsM���7:1�M���Wf�#�t�=�X�~r�o�ާ%/��C>s{H�©���͇��1|W�.�\�)�a&��S��ɩ�uS:�{�#��W��b?<G�u�3���W�����>]���[��z�7-W9G�\�K��1�% Ht4'N��\�Ƨ�	<J	PCp,?"�<A�9m�-oaT��Y�#���X�
�T��w^��#�|���f͙Q��4bJp�w� ~��m���,���Ʃ�1Et�ܱ��HDgd�_��s�3aD��j��6)�UFB�/����ك!Ɠ�S���[5C|�~���S�Ґqa�"v�n?L��7��uen�|;�����ӈ
v3�OI�<��k��o�8���M�ר2hܽ�N�{c!od��Fj�*�F9�;mKJD٠!$q�[E��$���V�!v5��I�"n��Zk��%�Z�rU���_�<r{@����4l���-޽����*��	5L
�����('��j�i������G�]R���tf߳�6:��P�<DK�k*��}g�4Q���D��pa!���.Yr*P>e�hDp��B�91o�1�yl���\Q-��O��O�ƿ��^i���KV`ML7<fP��j�)*���v
����97^D��!b]Ӏ����(�o%=у��G,.���kl(�)�-�CY�2ءT���e?_�C�l��D�c��}��Jx�U��}��H�q���h4M���x+k�r�`��5��j���D��L�vk���^��d����~p��`_YO�r��ݗ�UR�ї�WH~�>���a\�|,����y�)�_Ġ�[��B�ׯ�GIy&p���4���ծ6�,�Eh�}h����:w-���Q$�����OEM������!]�v>|V�jP
?Q���`����j����q�G�����k�[��U<{������6Ho���e�+]��7dA;$=�f&S�̀,�����oa�`�2-�F[w�b��s�w��z��W��D�hp�e�V*��z�N�T��D	��P4��a[�b~�l�w\�Ni��UI��C�[��9X)8,&�IA�:-��@�{+�> �s*sS��B���JX~o����7�&LGD��q&Ӎ�UȤ�sH����'F���VΞ����By0�%�&Y�AFc 	���M��Q/Ҡ�lX���t/�[�S_Һ�g�
�"#����1���b�-�����X���t�t�
������I�׵���͠��j�]~��7���I�?�LT�ɂ1�V��JY��j&���z��.�d�<m��R'j��#����L�lyX�/�U�+�1��f퓗p.�"9�_8���݌���L����&�+���m��^ԫu�]Y���
c?�N��
����TH�Q��;��������ě�{��`ܨ�-,��~�_��mc�D�����m��g��$���v�+"ʕ��/���~�C-ׯ�t�z
�Ma�U�t�FKև���ܾ��Y?��;���ɣ3�'�Q���Z��l|O�\/3L'n��4�Q� f�����>