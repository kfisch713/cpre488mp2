XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���m�Iy�g'>� H�k*���������}�~��� gE��'Df]�;ѿ�g��[��Ͷt;�E��r@�B�;�\��s1���Q�x��h=������Vl�.F�R��Z\�%[d�|t��s@��(k���ʠ��#3z�������^���.�n�s���ibX���}�:���Y�Tp*�@P�����\j���������Bm"�#J6��\�m{���1�.>��,���Slʪu�m���5���ՕL7@ny��Y��4לk~�����(ǃ�ʏ:�(��p�oD�y4J�xx�37�D�5e8� dR߀Ѩ���r�vm�#���)V�n3JO)��E�鄊���'S�8����D;�����Q�'t���4����[2�rD{�eү�ڧbw'��Z|���=���]p~:��}(���W�����-�W��d0m�K�l�/�C��ٱ���h�A�RV+o�z�m��q�OOF��J�"s��t=�;!�g����P�EJ�Q��,�������tۄ�E�nŶ�ʑ0R�I="^�W;����#�����6��������Ef� ���W۾��'֋y�ՠ�,�?'�,i}� -��3!��
�9���ǭ��rW��������.�o�{ߝ�)�ՄC؞��l���΂��ުߴ�ވֻ\�"J���9�U8�j?F�H\���8r�q�V�}S_����?1r�=�uP����Ʃ5�M7δ7	�-}%����d��`�M��3�<DXlxVHYEB    3b09     f80���cM.t3��!��:�=g�b��m׆1�Chnfd/HG��E(UdX��vj9������}|�A�Ye�ō�̙~>��`�e��ug��N�<�;u4VZ��w��y=.xD`y�I7e~�G�Z�}�ؗl�/���U���)��HT;�32��y���I��wy�t�?[���Θ;T���!�ԛÙ`�C�J�� >�>���ڕ.עJ%��W_�W�gA��ԥ(��MT�w��G�f���Q͓���#4/K�~i�z�awor�����[�z��Nu}�na<P�q��_��@����y44=�G�G�{��oZ��<�8&�8�qD�6�b��ŠBʓ?��d�2�s�bـc�c`eB���|V1�w���ڥgZHD�q���P���Y�H�C����lN����|8!���;�`���K�`�]����?���)�a�Ux���YRx�/�X�9�qn�I��<�z����@=�g�B�O͠.��*��Qޖd�����d�~ގ:�4��j݂i(�]��wM�h���#`ݐُZ,��w����$V��ǑTb�����a�T��ґlv�iO¤��cvd�>=�Bޣ8$��}[&AtU5n9���;����&1�O��aL�t	]r&��YK�{��_͛`��v��
�\$="��MG���}�� 8J(
��2�A�)�Zy�\���p��YO�z����F1�����\V\��L�{`M��l9�$�|(?��
��Ї�zZS��{��F��~��;�Ϻ�!|�6H�^L2�;�����Q��/���G�W"
��l �H��
��{[�x�Ӿ�J�����¾���8s�Dlu��8tt�ʰ�x�ۻi�h�hB�"7&���XkQt�Ib�ນD���\�+�Ǉhfﺭ�;�h�:-]׶����$�W�!��MӶ��ӡ5�[J˨I�?�ֱ���˨y�{�K��{9��]��z�*������:�ɓ�ه8|�}�S.S�5�w�D���y�  ��шB�w�m�J�� �R�zɥ�I�[U*51ַ[r> u��]��^s�t9���oM�z>�Ô|��	�ծ�H�M=�`�gU ��|����-�>�-@����,�5'gݖP�|��?��E��{RV33�L����#j��t�P��\�v�CDDO�T�jm���,�,��Hdҟ���!l�
��!Y���p<Xr�"�ot_8?4��P���Q�M6-���Øj��h�Y��U�w��lI�RP����+`����@xDo׋K?�Wv���K�ۑ���%�]���r#�\���S��T�=�qd7��!�J�*�����fU3B~�������&�^��x��Ѡq��a��*ض"��b�����r���@�K�Z?卩�[K	�|�RHhCZ�D��E-<~g�zy�<����{c��'a�
'n{���MQ�4����M�d% ՛|^z,9�`ԩ*}Vђ\��0(!o)��%�gdC���u�Z��CE�w����Y�w�����1�2��+���%��{z7c/�8yט�C�`��;�dXB�G)8�}�<W{��;D�?F��=P��T�0�~rF2�|�)�]i�u~�����H2��]:�IM �����#!��/+��
�I��ܧ8fb�6|(��/i���ϖ�|�Z�"#CIҦ6�΢���A�0�-/��A/�����,�!f��3�����(V˽g(�E]9��U�P#���XZF�A�8�dl��\�+��R�|��_;�D�[R�y�$�uH�.i5�J��$&+UU9)@	*Ă�j9;-�p�w�
.a�^�0_{�X���#�\F�h,�o�5 �yy�����w�_>tG�0�p�v�<r7�6��8�> fn^h\�wV�Rt��A^7.*��_<�k^'AL���A���1ÏUk'���U!���\J�7L��<�����除l���CI�@��A(����,ay͂�4�ɏ'C����t�Z0N��
*���`������)5���c/��o��	��m���v�h*u����*�{	�4j�ˎ�J�w&����oj�ͣ�y������}r��8`��f�V���g/�k��2?�Og�p�J�y���4	������ƹ�{mp��&e�eD�Np���K�9�a�I�ά���ܧ�C�bQ��yn�	��iM�<91�y����P���l�?(G�LD	�x	5Q�`is�h����$�ѷ��6�t%��Gn�ZF�ɭh�<2���Ї��f�F��&z���3*N���OI�>&0�p��fPz/��(��Upxy2z��Øz����>u�ݙDH�_�A�^��_4\�ωY8HХS��8v[�b4�
J5�q��,bF��`�3tB>�L�}�����ʑ�E\����ў`h��Y郞~����"�ξƮ�B>i��>x�UM���ƛa�.ƹl�����3�`?%�Pi����r�^���}��r����dPh@�qP|���B�o�/KHt�kŤ���6.t��������1�_N7��S�P��L�7��=d��#U�����h3ə�oϦ$=���l2H6��7� �h�?R�ai*��P����J2�ΥPs2��M��|)�|�@����%���F�u���C��lΡ��(��]2��.8�<}��y���U���ӄ�Oy�Q�t w�{!���Ï
b[�Tc�(HO5X��s�km�W����%�A��sY"��`��F}���ĵ����h��:	�,�3�~���gq&���AeC�R�{����g����jNt���䇂y�tM��;̾Kj�:�ș] �S	6��ݨC�֓û����C�r�.�A{�w��J,�;�(�ܮ/���)	�c���Z�-2<H�XVNǓ��'�Rޓ��ʒ�Q����׏VZ%�t0��1�#7����.�#�1C��۱�O�H�ԓ��������XȀ�u%��u�T7_D�?�m��F��S�ǰ �>���o	��g��u�\�x9~����+��ec({��?��Q����k��=���7�}�]��Q~ˬ2���:?T� a��
zۤ�D���	W
�Ǣ?��󣤑�d���n�d;��A[�h����tI_����{]��Z).��� ��|;��Nv���`8��Y�nPF�yo_r��\�+4i+1ܫ��fo�dh�Q�A�nC��}�47d���<�'�4�0:v��o�_2Z0�T*�5����
�B EI��^�4.�Śde�0W��	�)&=��(��@Qdvf<�{"�f�>�yQ����"j_�-;�:��za����Hf�q���.�@|��<�K�].Z�u}��
ڜ4����Q\�d�EW_ S�jƬ��PɎh�/ ���B=Ir�U���nW8��ۧ��UC��ΐ^�&��V)�}��ן�J:��Q�`�.��L��nIR���*���@�G�$�a���Z�<�<�*��]v�`����ۊՑ�S��V+g��Q����L���̗�y����f}fr�J��\D<"��P�ժi����l���QQ�N�����}&��h<���]�[�F���KG�m"}��dd_<��c�y��ZM��U �|����2㾨3�����$��'P��x��`�rA�c4�|&����2�����n�yIb�|S���
�Ј??�gX}l�_1�5��O�<�'�$��6�W=��6|� �"�gF��_$-nc4T4d�jJ������o=#�y��7��E\fw�xoP:�>��x�����������!B��<���˓CXbs�e�%�?��0w���ķȃjx���#&�P�����a7\i�~j��U�N��t�R��U����AФ�=&�91�lP|z2�{_�Q��E��|]-��