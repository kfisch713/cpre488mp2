XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �\��_��x��Kl�׮_q���E�u&��!h�3�K���~q�z\×���l����*�>�G�Yt&ԛ'�8�sf��If���;���LԶ��O[�K.��d�K���$TS�R9o~�]��(����W�-��Vl�R�z�2����i��eb�|.����͟������P Tu���"*�:�6�	عE~#�,�֎�U	�c#"�"W^T�/	�.�G�K�˅-�@.>��o�5�����A[�GA� `	F�3ީ���&�+*/=q��Q����A��y#�x��i���~4d��Z��B�X�d?2�;{8�^�Kw�*�. �ó%��.7}J����+o��
��|��I9v=��(�j͔O�JJ��]r�S��5�,~��π8%�տ��z8��U7�A���e�<��w��ޕ8�P&ѫ
+�x�0��i0��=�\^��]pP�-SP��p����[ػ��?٫�����s�č<�2������Ԑ'ϊ$��l/�9}�k��"ެI4��;U�U���2Q��2�-,v?�%�_�T����a��f��ͨH���F���7�%�`j���TZ�o_ޒv�E5�l#�s����(�C
f���,��^�*�aN+�w�JrT9����`ݚ�ծ���`�P�_�l�fV������j9n�| ��Ґ������oCxp��b.��B�9Z��I�f-�$�%�>�����D�����l��O��K��E���@��\��Xgʛ9a�rv*���!�XlxVHYEB    82c3    1970;�j.��O�;@��t��4������Ҷ3�
/X��&��УnC{���Jd��R_�E�[��,N��~?�sD�t~v� �ӏ�VFmu�u�փ��,ޤ���-��2Łj�s�͉����(u����|4�g�|�|���l��hH��O3���j����m5ﰆ �
*`�@�}���O�|`��>_
k���\�k&��p��"�i�����1�h;ĵ�k*
�_<3�v���2-u�A�c��ۇ��6l!j�'í����+Arj1͒�i��2�r��(�a���PJ�+ڥD2��$�$�HY-�e���-ԫx�����0ۨ�0��Me�LpR� p�@�n�>�Ɇ�B���7J��Thl���?�@7�J���j��-S7Ѳļ�W����)�1��\f0Ù������Wu/Mb��k��Ջ?���Z��2�@���4ԢR��%�4�0�;���!ZV[���Aq�?��{����'�&�g�(ODV�Ov�(߇�j3V�]����*���!�F�0,.��tp��c�9s���n#T�?� j�s�E���Ru>�~�1)�2�	��C&D[�i�5:�߁�1�aѢ��Y1��:U�r'�;�����Bsf�V_���ܦ�?x&�=�hf���Ħ��Y8"~�VG�9�u��*�5o�s�	�����[.��{���P����H㑭A���W���(��L&�;Adh�S����څ�5����r<K��� ]��Ώ#x�d{��_��*�����V�q��A�J�0O�ȡt1��ț���s�:�Nh�tH4;A4p��^n����_�r[��xd�8�y���^S����e�).��UѮ�)�F�UyE�7և"�=�������Y_
М)3vO�{IE�)�bmڔ��w�V bFa,`F �{~O��u�z�F�:`>ߐv�'�ҖG�;�Q��Z�#U+A�ȶM���Iw`%˽JqM�Dv��=����y�{�w�_�X9㫥_<�AX����+�k�/��w���ǿŦ&���o�ŒH�㧷�'Uȉ�ɕPK	��mi�z��^#����x=@͜�v���;3�x�BB0�7�ɦ^�i7L_�rw�n�O�?�5�.�1>VR9��߈�Å9唪P��c�Z��(��F�a�D�5<v�A�ǥ��,cǾ�i�^i��!lJ$>��N�֥ "|�Zj�V:|�2Ö'�׹���?�6���z�h��0���b���	�`+�G ���H��h�쨊-*w��#�I �T��2�� �fY��ė��Avd�t�k�J�{W�	�vw��]�=�˄���C2#�G����?s+�a�7��CG�{2��x�Z��Î!�']�Ibr��Wא�HV�µ����Ti����'�x��R�>"�[�5ii��H������,�3��6&>s�߳���a�W�T�*�f�J�y��bc@������+p�]Q��^�i��+�C�ꉝ
p�w�C0���G�&K�&%�c	��f��f`���Vԏh�6�Y�i��p��<���Y�����_���,��g��?<��l���t$n�9
���|y�_6�<�F����pl��CF�x&�+�Y��;ws?� x�`}�y�B٤߼�H����/on6VT5�n�eɻ���^�Y���>�VN�zܒ"������轂	�;�u�Er0ji����(���d�#��o(�`�fT����yH��xV�J'S��5��nRn	���� i�n�Cic�hO)�Z1��l�2Fa�8'?F�֯m�`�h]o�1�y�[�'��W9���%�[���6f��O���o��{ ,�`ӆ��:b�ݟf�g�ѓ��Ҟ�4eS��c�^���Sz�r.xj���Eκ�d
!r$9ѽ���H��H�Z� �)xs5�Œ����=!�@� �+����b�9���8
��d�c�'٬y6��_����E�`D�j���R��f����3���k��e���5�?A�:��3����t�x^����w�o�C���-4�>I�r��](
оsi�e	t��&2R�t�� g�ED�����b��jg=+��m}Z*��/b�"yb�_���1L�$M�U��Ͻ	;)��� 3y�� �['��f�e/^�J�TH��-�Z,���r�n�$8��1~�䝇�q�n��{�;�<�3��JY��4GR!"z�[C���R��`�R����Vy��^�Ɂ�j�P���`�g7��i2j�f`nw'����Zn��W_��j�������G#U��
([ŷ�Thd�F�^nyz���p4XՓ�>�t�[���EL0t8o	�U	s��L�!4EZ�ќ�������۠NC&�Zk�#�	N:W�� 7��o�	T�Y�Rn������K��W�]�c����$w�L٥�q�e��P��F�9�w�$w�ʚ� 3B�!�PO��Ih�H��	Ȝ�k����x�wP��'Sy�7{�'�""��b�ȝ���:2z��Qs��m���u���G喁0�=Τ��Jedg�s��z��E��Z	~�t<�ւ�E-*�<m�y U���C��^%�{`����$���-�N���5E�zy�1��f��3�ӥ���*�u�xD~�1�B����Gc[ �u�j�$�l}�<;��:lo�%9b�.��/8y���>�a6i3�g�i���ݵH-t*l*���950}P�)�N#��h��&?�>4�N�����w�>}5���_�Л�6��/��!Eb���]�E�O�!AcU�G9r�������Q��J��T7��d*����Nc���K8������rE�\O@a�"ϥr��ژ�T�ީ}�yw C�1	�_f��8�w
&�ˋ���������طؑ�1yK�����q��A�{��M��xx�>�vB�A6n?��?��[s brT�	͓��&���3�Y^@��&��� ��*m��g��ݳ�J��7ҍ'=�5��� �����`��1@��ton�����x+M>�4iM`�֠��6[����b�v/�hֱ��3)f��u}�OI�����<��E���?��>��z�6�b�q󻓣#�q2��6�8Vð��U���� ��֭��`�ĕX���[8��q�s"M�ua���J��P(��W��2���/ל,��j�rl��WyZ`�hp2��O����C+Ƙ��c��<	URNDP����6��d��+N&AЬr}�	x�Hl#?�)3YM�����Y	�W��:`�m�sh��'��R<�.�Ι+!��Ă��¹h9�D�����)����"�`;8�>V���Q2�r+U9 cZ��˒�_�Ǻ%�yӸ޾��G��IYR��0��[C���4k�r/�4���{�f�u.=R�Ԯ�S�*j}7�#�osg iyC�0]f�5�!�(0(L�8�h.}yr;:L��e�P3:��;!~o�ś�y�G�8 �����5������8$�y$R��#���v����l��>V�S��7w����п�e��!D���A�̹5�]�Ae������G�m����9����ܯm���-䉋9�`��C%?1 �S�Ję����F��lm5n
r͊(��3l>M�˓�x���`�	'�&_

��Pļ[�^�/�qQ��.����cr�q��Aӎ������XjR;ٕ݅�Bٚ��v�?��5��Jڜ,&�_Q�����1�`��lz8�z*�V�;�:d�ش����}}sm���������̧P@=`�J?���w�;G���V���Q`|6U0_��V��H9��	�d����g�P���g������W�Avg��[�м�Apڊ����	7�e�C��S������R��鏌��SN�y�,�E�ܔ��Y4Om�FI��'����p*I�C�Yφ�M5�ٹ�p%�j�!l�([��r���Sh?�G�!�6��u����.T^�ԗ��d�ւ��8�\m�ז��r�/ôۉ-�}㏐���_)B%�I�^��;6�R;��fd��}���h�z}�㘈~�H����^4��,��{���h�}jl�ZA�	")nK�[�ҿn���@�/�szs_T���ʘ)w"m�&��q��������;�:6���5�%��sǄy�
���7y�Q�6�W��5'73u���A?l����R�6���W��%�����.&_��ɛaIwezM�$�A/�!6E~����rOhΰHOlL���[)��8�7�={r��Y	wȑ���S,��� �gRMLu���%�a(�&��bM��(��ƨ1p��_��&Pb�N�'�)�D�a%"i�go��~]���e���+*�z�R�g�����Y��.�8���tg��9% ��-�4����1�M4��{�ƿ22��*0s�Ge&�>F��˶��u��/�;R3P�>n�6cˊwQ9���������O_)�t/�"�,D�/�D�>KW褬���'�f1f�ı��|�+e��~�����6��6�Di�J��f7[��%����
{gߵ��8ގ*D�f��L��
6�f��e�;>������`eùԈ����Y�1�2V�������~�w�	 .%k�lGM����8M��@����k��q���N���8}�|XmO��}ǭ��zY�w��v�߃�0���6�2�����)F�ѱ��ZM�M�ǠC)�t��ZCK{w�U)DG�w�d��m����9ɿ]V�=�5/	����e�p�
� ��t�/��͝4��l4F�h/�޲�����jR�`Z�ky�p�F����n�y��qԟ�݅�\HH|�D@z�-�����-p��&mS��y�B��B<��E�?y���t� �$j�bV���A	NL�!�G�KY6e���� n��U�l�Z)�3��>Eq������ޘ�`����e��'�,,�Ye\�j/��;�N%*�t�E÷*�-^s�1Q�H�B�_N5a�+@Pʅ��Fox>*�(7��t�����,�s����5l�[�=�1��؅]������#�I��Ô�k~����I
\zH52J����ׁ/�L���p���~Vg`{���E +�_�{ ��N46(���*�R?f# ���[��W@�3n}�,�Q8�9����
q�U����b�2QS>4O�i���乨/��b�܄=-��޽�f�?vp{�u:���!��n����AĖC��B�lT�S(ta�BFy-tFi%��<�وeDf�r��ޖ^ZZ�%z��=��։)j*iO����c���,1��) �Ō��m��ej��2��n�ƭC�SG�1��!}h˟��x
�!�4����T�a�`�z�_��ZϪ�dx��A햳�?��mv��G놠p�r�}�>*���19����b��UH�;2>���d�̀�'Ivj�Q6�̂�W��>>n7�n�G�I���5��Qj�X��6M��@��0sWx*+"q�X#��Ba;N�28>ׇ?i�bը���]�Ol�L>�_��&8�xD)=&B�5��n�M�Ke=���t�5~�����Ft��G��=¶13�d�;CGeIt�B�'���f�M�
���}J���rZvC��H�&��bb3Xd��P#��	�;�Gr�����\�;��Ac�QP�.\&ρ��m�	��s�������=6�W��ǈ9Cw@iߘO.��^!l�i�-#"[�#`[�m{�%A�T���H�Αi.a,��!U���շ�Ξ{��t���Dדʢ�b@UlL���U�.��ts�ޞ7�}���Hs$��\���R�(�K�x���Ck���}#��q�eat}��B�����I�������J02rqM�7C�U�j����~+=@ģm���J)8k�4��q��Շ Pצ�z�l�#x
~<I��Z.>�໲�1��3P���uh3s�Ͽ���V�J+���i3�����=*�qhDf����K�J����d���1�a�m�����g�b�e�-"�!V�(�:X�<�O�auE�@}_��/���*�{m9>o�6˱]@�qx��;�y��Q*X�42ٛS�Cb���.�J��%�n� V����v������\�Bj��kR}��#����,�r��u��|���,����^VyrQ�C1*U��X�x)�a��
�Q�\���;���,�8�c�b�?}���L� z52�:.>�%��U��gQ��T c�E�	%2 \���d��ӹ��+B�,��w�$b-�=	���m��$`zfP*]��xd�P����Ϯ��$������a��=M�5F:s�W����#5��{�3�	Y�������Ϗ���k����/�
B&2��V�>�a��G�������G�r$�7�8�I�ץw4����L�GG�j���i�ΫG��6Wy�Ł:1K�w5Nxg	lx���9#@spR�nH{?