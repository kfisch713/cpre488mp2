XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����!;�F�p}�nt-Ƅ��SY[�7��B-S���K=�ӅM��q���"d͠���`�]�ȧ��k/��MBQ��s�F��k�2Z�y~�*��y��H�{��j���zx��3���,S$��m[���=L�AY��²��R��4Ms��F��!ǯ�`�N���P�@@'+�p̸$�)��姫�(��Cԛ��.Jɯ)o+>�1��^L�%�ê/?�Dx4�.`r��Wf׃g�>k�wrl;At��n}Ӝ���IF@�G%��Ɋ4:���/�s�����W5���bE�(�k��u�K�_����N��*9sc����9p� k�}�i����P�<�F�~R��8+�_!~�̼��򧿡�*�H)��6�Łx��$�	�D=E��P| cy��뫀t}ʠ�IN*ņ���xR�Bc,��ϒȨwZ�V&��I����Za�C|ަI��Y�r�b�r͉=]u�M��g�C�rb��["m�-e�Vp�9ךR�������W4�|����L�]:t�_�Tص�n�#d��k41{my��<�������b{�>ܸ���ږ�	���$u��Ʀ>]N�~w�����o�s h�����4���	�+U��2庎0\���S�[��m�M������kZj�g�� ϴl~X��i5��RM�;��/���
@�J)�w��7�¼=�#�ji�U �V��Y`}I�Bc��_��g���X����qM�d�}B�%����<������[��+aD�<XlxVHYEB    76a7    17c0F�t�"�W�R��ڻR�]�u9�� ���.BC��\+�~�V#7ޙ)X~/�U�ɇY�F�R}���"
��[�a�z�L��kK_�Ą�_J���F�e���-.Rڣ�`�F�i؄���ot��	~h��EG�&�/��z;ݲ�TΡ��j!�t����,�	����<�Ҽ�-����u4"��N���ȭ;f/$F4��5;JL��3o<�𶩉1���Y=����yFp����!���F̬Gw�.�lk:�۴▂ρ.�������\���
@�~A�!��ӧa@$���X��8
 |`9�t��Q�F��V�Ȭ��D��<�S���#,�a��0��m���b�#�a���	�����[b]��yQr�"��:♕��ĆK��iz9���M��Uu�q�X�����<0' ����5雝�&��0�1o�[+@X���gu�� ?��q���)�5Bא��#���*U���/Ĩ�xR.R���L��+sJ���5�6q���2W0��m,�Β����b��){�$%"=�ԝuP"��{m�H���.��M�ʲ�מ.�Q^�}sAҖ��:Z�7'���B��m��� �mZ�^�]k֦��`��Z��$��LEL����7n�������Y�ª��.�&�,a��{�MSl�)g�oo��������ZJ�Cd�G�U��e=7��|:ŖRzP�0�;�A�V_�Y]�2%֞X� H{%89ٞh��+},r�����o�Hag��N�/C��QߤF*�@w�F��°�OJo�5Q�֠S��,�V\�x4�*]ꆷrY%��� Ư��2\2`�{��V��l����0Aw{l�b��Gi��u��x���
�W��g��q!X�a&1�\��d�������2ݔ��Y�=?�:�i�e6����?c6�	^'(���Q^O�]$F��Qpl���8*�	��E���W�K̴��豖��0�m�Â+Kp��@�:o���rl�?�����n��=�$��;רr��L?���bk�r�g��W喹m_k#6�X%��489Ĉ竆�lTqo�e`8|[����%?R���zC�E!^��a�0��t���,.~-�M�_�ۍ����k��~-LG,��2.gl�X��-B�� H(�A�2�M_p�Q�_��ޖ�����L���o-+9��Cg�*��k�!��8�<�D�r���C�q�rD4/~��?���w̦�	'S�����IdǜF����E��4��ɩ��4��B��$F�x;��]�����t�a{a���0�D��t�Jk?��H���j:�i��*�����HQ�,��!P���7��!��$���Mm�ߥٕ���DwG�΄�Z�ϑ�PF�bY;(h��A��\�������Ҵ�:"Y%~���?rF��\��J�k�������&�a�|�s�$c����S�}C=�/UX�N��に���0��˽��W՟�0����8Q�P��uI*���	��k�~�� :����F��v�:��C�8NTܜ;�^�):RJm�s�%n�'�4-����a�ސ�6�p�-Lll�����YG/��Y���R.��-]"��8�+d���n�,׃{12%� [o9�f/p�A٫�t$Ű��!���ʼ��H% g���KE�q�f6NW���G�C����
�G��<U=���e���f=&���/���3KC�N��f�!0�5B6���t�~�F��%"!Z����Bv��]�S��uOv��V��9���疳^&%}n:~ �ք.��5ۓ�F_�$������,w�h� ow-/e�����.��Un�o�_U!9�Nnx<�>��5�
�Gq8#����H���2�T�]�ۈ�Jɾ���1�䤁b�B϶�\�4Q���1y��D���D�)p�eǶ3k��$��Ȝ+�r������=,�4ъ�}����mMec\�	7 �\t�\5���o�����r�B!Z%߳�;���ݔ^_���Y���$�D�C��Y5�C"r3���I�+�=�d��Ũ"8y��a���E�8d&G'�v4g��GNJ1�TS�{�Ĳ�ؐ9�3��rU:��3�k8ܵ5k3U!���� ��F��4��+�������\�5�1�N K��eM9K�S!�vV�c�Dh":���e��筅\�fy�0���&<Wo_�B(0�כ���\����P���5��$�i��'���Ik�yb���!��`a����5�0�-2/��W@W8������ �ذE�����}��L{C,?4�<<���Գp+V���{2W���`�=�A��_rK 
�o�_���0^A?���q�tsU��p6ۆ��}L�Z���h���m��!;%	�'�Bñ��dt�;G�R+��=�E����ǩx7��d�V� �4򘄠k��ᶲA��=}G�t��82���1v�uRظd;1�a1�n��3%��$H�R��X�X�=����p���3�/YM���㹇/DC|�tYAq�ˎ���R~2�B�۸!5,Z���S���]-�.��V�Ҟ"_}sݯ�2@xR���ⶫ�
էԹ�g���o?p���6l�C�2խ��P�"~��Ⱥ�A�6K]�3£��&��3��7I�[/���(�s2O`�=��=�Bt҇{�:I��o4�Zm	l+�0P�%<� �sZRp���(���������Ο�/���6�eںY$�]�:��OebO
"�te�ǫp��R���.M ���:Yf�֝���6�*�0�J�ެBW����I!8�л�\��d�ޱ���2����6�2�mh��#����ۃ�����N	#���	;a�[ǽ�iS3\����inS�z��N��r�aOw[|3ClŜ�Ϗ��Ϡ+
�W�-��d6j�|&���F̟�<�r��۠�8ŝ%A.��s6$�2�hz�ךӂP?+�E�����JJ�ȼ`}.��s �e>�mthW��N���
�O&�r�;�>`E� q=],d�ȧ�L�����6�
���=��M&7�������)ՎYm�7ɗpę�����b2iұ�	�D`G	`�#)0�}�q���U����E
o��>4h1ɠ�ݦ/�P�"��H�~xPb� �)�5��d�ٟ>9'Ͽۊ�$xH�o�/\���6��3��U�s��[�z�����>�AE�~W����L�@<��tQ�^�2�����d���������~އ|4E��%}rKZ~�00Q���A )��1eo��B�1���Q����C�U*Y��(��Z̞&�	��J��=�i���Ŝ��4��?��v�ś�-��F��8�=��F��9��Y�0U9��,�����-���Y6̨��:��pӋ�+�?[8�7Cή+><J�$��3��2c�>��Ӷ~�x
���5=��A��C���`RCP�$3웓��Z$�Z���(�9F������rO����#���c駘y�B�/�����̫���<��k��+�����뎣V7���zDd��{G�����j��`S��Y�l���2��������#���}-6n���ɱ���q�
�M�M8`�|#�CX�������sj�%~|��EG�-`�D�;��XBk�v? d�`��E�8S �����ʤ1�E��/G�{iĩ�������]��k|١�wv09���A�к$E��&�,I�^����F���>[*�� 1�� �0V�/��V�������V*�{1dx��S�Tx�#��Ep�;0����)ٷ�V��x�������c�wAlJQF�?����6�,l�����gO�fDG�7��^\�$���7E�;۞R	����/g��H�6�l�bS�b�^!�C�u�^=3#��H��2%��Ő���c�׽��Zb���Z�	v/V��/�iCS����R�K[f�9zh�7!.�k����\�Ź�f�x�{�v]�D�?���}[e{%���ݚ!���,6P6	���KBZ�pY�$a�:��]�X��8�������Z�A�|���@�e]����X�ɉb��b�P�	(
��qd	]�ſ[��y�p7�'�*4[
���Ԉ�����y�v_��1�f:��CnH;�BI�v�S�0� ���E�/��3�/���i�9vڇ���5�/��A��z��*�an}��A�hg����@w
!�n������`F0bEm�l���sC�\2~���M��vCwa����z�ކ7�l�6�꛻���6��c�!�q>�26�G�������*ceBss��m	�K=G%�/*N�䵰+��u0F��Eu$�������Gp �0�P��3HM �|j,NB�"���jx[����m7�&K��b�IQ{PI[��Z��Ep��V��b6�|��ax�����V7�V�1��e��!�
�'���`�jP�Yg���V]:��W� d��j�=`W��L��I�k~��19�J��9���*w������@J��ͷ���$�+��-��|oWॶ`�O��ٵ̛պ�bd���R�)Kf~>BZMr�P �<2��s�6����N�#fS�}��;[&�aC"A��&�.�S�&L�w�GE����-՟e�fِ<���q���K�����6Z�=T�M(#��H0�����6��~#\�m��$2�֞�w��+��V��E��&��sc��n3���>m��s��1u_��8�k	�Y�oa9tc��cc:�ィ�I�)�?��d����w΋�ML ���e�RaI4Z���x1Ǎ~��4v�� _�8Vq
�C
Zfܝ F@cӌ�'�P�T��,�t���ϕ���A�,�k�;6Y��j�����sW� �<Z�� ����"����㔸�s �X��G$��	�7X�f�0E"Ml�>�^���I*ܷR�<�������q_�zx��J���
I*70��W�'�X&� Mt}q�4�c&8^cŒ������9KiM���vǣL9�6�b��ߣY�*T�NP���p�=g��(����9@2�kj�i�]�SWbH���?}ñ71�hrF[&���'�64���u�L�,1R��ٽ�=��K8E�Iy���ev�NtUb uE_�ޅv�^�9j����c��9)�헸c*������=��)sf�������+C���M��5r�ʊ�>yѰ�fl"䦳
S'�m���P��ս� �ॖ4bJt�5rOg�/��a�`�://�����
�|!�6!%f_#��QT\oIq-G<n� ��%��X}7ω��X�n��c��y�i�&l�fC����K���ѵ4I9a@`#��ѡ4f���3J���ʢf���g8���RI�u��h�3	�_K4�~B鷶p]�0r�Օ>�"�ڛB`�f"'���X��*�;͸���������'�����|j��=���z�����ѯ"�ia{C!�g��܊�z�%��Woo�Y뢟� z	6��=T�n}�~��`�gD�mQ��>al8����CVy��0�wv�#o��?��@�'�;�%��SK���	���c0\"ޗ&����ת5+8�Œ�Շ�c%���uMB�<�i�ڔflD(檀�~� �z���[���e�r�:]��77��I���������G��mNy*1��MN���Ł��F�v�������;��~�O�Z�r�1a17�Y�t:�`���ԭ�q��Z�O-��=FN�z�a�7��I����+U��q����7b�6�)����?Q�9�D��nP���D�&�4[���
I����חe�V��a����h#�ڒ	������P܀���ѡ�O�Ŕ��P��(L�0��@�éq�}�@�Z-p�|��U-|Ys����H<��,]��H��j�	o���\)�(�%4���5bU׈�Տ^'5�[ ޟt�=��*j �}�m��#c	�k}�}�b������b�u��i=.��J?�fo�U��Ai�m}Ն�*���M9!@�h�ғ_u.	�X�eT�0���l�p��`�-g}L�I�/6����WN���&1��o�h�^�