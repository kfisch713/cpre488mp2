XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Evn�4��(~ы��8*f����b��������>���G��Gt�61U�S��s;��c5Ѓ�m&1q
� �P�Xs�!��Z��q0���% ��.�䦿�x��� ��?���"�vL̛���LrC5_ߧQ�������j~c���J C��Il�礪b}�+W�A	1����(,`]u =�a͘�pØ%Pe��&��5I�G�8�֓k��Y�7/X��W0{9��eF �~0=�ZA����P���gH����)�V�T��7jU>���3�/L���R o��R�+�ӊ��uѴs���M�!�4� ��%I�_W��$x�/��l<ɚ�л
����\6w\�D�u����=w�%���!�c�g���P��{;�i�0	 e������+_����� ���Cچ{��Y�ܶ�'l#�)[�'`�Ρ&L�=K"�m������bf�y��w��L�睒E������҂M���m�}����y����Xf�Y�TWR�}�.G��"c5���]u�@�cX��3�>��4�ŏv�>���u�;g�x�%�����#�_E�A�dA&�R1�h!D��S��j�
a�@w���K Bv�9�?�B��`uյF�T�e0�����$�.��l�jJ�PD�f������(�A�G*�GS�R$�������kM�K�Fy�շ�T?�9M�)�����}ʕˈ@E��UV���jϠ�������ZH!�0��q�D��X���XlxVHYEB    5d54    14e0<^u�}���{�C�t���߶�U��=�2q�B^�j�G]؂���H2Ϧ�-
�,�dL�
��r���a����4����a�Z�D���l5NgVz��ǹ�|���^U��k��7��Aw�M<Rc����
Ax��=��&�h-�
�S�=S��wt�Jb2��x%#�*�Y�y�_���$C�x9���)?��b�#`�J`-�C�EcL�d�A:�0pe��2�عm�RS���J�p}���R�\�j5h��S�̕�ݪ�
�,A�CW��	�����ghLb���<
��̪�ȇ��6��^�gA�СG��'R���\tW]�x�K��}
˝ܾ%�^pgp?XW�69�k�ZYb����iO�<���� ��_	�'6�����7.�
4om����Oi�&x��l��Ь��g�A�Q��Y�(�T1�7�*9��m��Hv�h{�U�X*Q�-��\���R��nH~)bR���4���[W"l��c=UXx��'�˾����y�.���wlz��L�����_@5:J�!2,G�'OqT���v6u��w4�����]gY�v.�����w#�Y�)��.��N�u�S�l;-LH�~��$�T5�`!�:LH����D�b��쀥��z*޹���<]`���O3` �:I�$y�'���׫M>�.�K�i�j͠oք����a���fܢB)��Eo���j��4j����',�N�z�t�;�C����;�	hDC��R�P��ޡ|Dw�M���nF���>v���*�|hc��8��Jl+M�\1!�:oT�t)y�� �us�(gI*ۮ��������"ӳ��l��	G�$9�*1�S��\w<ݞ>�	�4�SZ�/�U���rN��k���lf��\J�K27���W~�A,O������}_��<�P�����=��h!%�T
[���8p)��[7�����^V%O��: �9�y�6" 94������r��	��{;-�C��}xe�2b�[c,���Ƒ�C��/��I�Wf�	
{Є᯺��VשTp?~���|��}N��-�&��4�M�Ҝs5ȹ�[8n��P
4��ߣ�B���B�US�E�0�0����+K���@T����[�­]�Z"ڍ`}69"��dl]�;�H\15�X!��GJxyŮ�F��3cK���j��٣��_�%��/�fSR�+���D��vG��̿
�Pi`�5�۱r�����4����/���B��9�r�@u���qL E����H:(B�nkÂmm����@�kf��}�0<��w���\�����0��0�k+"���m�=߸��?t��~=̧��}���#�D�L@ն?_�|�A�(��D׽ 09שuQG�'x,�W}/�)�j�|7f!|����X�����A(���h3�z%�A����a��O]`1Nj3,�3��D�|u9e}���ٗ��l~>>�\-$�<�X^���0`��9O����ۍ��sG&9�k�B���<��A�E�����ms_��)f�O&����1[����kcˏR��\&��N�����y J��[s�A�2�/�zK�S�#�A��z�������/l
�O�ѯ���'�f,�gXKk�1x��q􋮙-'[�6�b���X�Ӹ�w&�2��
���Q��+�tL�-�܉�'�V�!�J'�lp�iڍ|/�zȂZෞǡ�XX�-���i�Z,��m��J�����3)��$D��o��HxqD��; �Ƨ�"�o�ՂQK#)K��Fc�i�s��(f"�\hh�� #u]�ڢ!0�o!��dӫ�R�o���g1g���9�Vhr$�K�/�QP��Q�aq�a|e�Θt��G��@ 2�v:��_j�U�?�I��d���f1��;�>f�/K�f� ^�As�^�&>ߜe��a*\F4`7Y�ɡ����n T���(�΄�2����j�N@kخ�G8
J]>��u{ֺ|
�F]6{�����x�V��a1�9����%�0���R�FXM��������j9 /����X�t��8^DM҂����q�Nj�e��'�/6T�0v��e�_��8���C+~��v�]�\V��tnZ��}�c4a���CC����.L5>��ߑ��ϥⰷ[<&�O堨��"*�AC��Q⠢����=�wB�N'�����fo�-^}��=C��ņ��Ӂf�|�v��89nx�J,f�����5��YL7@�O�\Û]c]�Ip/��$���,ENO	����ȢDb�eML|6A���~h%���䧘�\���BJZ�e3�D�e�En�]teK����hޘu	�g�"wRS��m��6�EG3K��ke,_�����_���c1�D�^}��K�Y��P��B�����>I��D��K6��Ap�pBPš��aí�5T����T�����7��A�R�{dý���%Lʱ!P�/���?�J�ol_�T��~0>���1����6��A�Գ�מڌ�l��[B3,\�)B�xt�,P"�<:�r)��<�}���xk���
n�t��V����}@[��f?���!�Bg��E�g���U�C"�L�tVַo������~��yu�d�dPsM1
=r�+Ta�����5�퐓�N	��,�&f�
�K��k�K�hTZ1�$u���`([}s.v����g2�d�_�N\�n�1��X�z��B�wd8с�2��k�8�0/��/h@%Cf>�>���C)�����J�Ӱ�uaH^Ys|"����+�� ��}b�G��@�*�K���h"�m������'����G5��K̤>4��O
PЬf��XV����75�8�.�!�H|	<ي�R_S�(X��gm�����N���:2Wm��ջ��߹�J%H��]~q���,9��d�='�1�i�	�Ss�Br'�����,��P��oNP���e��tB�)������(np�AVᰛ�"���;Ѽ���)e�B2I�O���;��QX^�y㴊{e�S�6��u��8%k+1�����8J=�"�!OV|��__�%~��k�f���Y�ݺ�z���f�t�H�E]��7$�d�FU#�r(ȃ ��I=��-��֪ ��r�%��E 3�e̸v��b6�ᗹ�e����vlz�&�g�.+d�^]�FѨm�0�c�w�1o=0�0����{�`j�۝R��)a�7т@�3�Y=��O�/K��_V���N���6��S��X>iM�Ш��R���Q��.Ty��]d+l;�M,�Q�3��G&p�4�4���$_h�L�|Q�ʬ>٘����-D�;�K1�����o�j�x��p�^)K!���8?ւ���'9_��ݸ���63���'6>;r��%�iAl�H�,ȼն��s��ơ7�/şd��9~�S�\͆��G�%y
��q�]��P�~�nG����]�Z%��P����4S	�\���9p��7u�̽��A��#�Xȑ�¢${��%�S�~��>X���J�1S �Lv��z���$_��&-�����`�:�ᵱ
`�
�(������g��2�mE�铱�������x�T���>�,z����&� ���lGJxt��!�u�������C�,���2\N��tϩTB�:xy�5y��lvl�5��aw&�m�y<�N�����G���A����<�C��I��<��ns/���%A|3K��2�\i�L�jc�	P8/W%�Z�"J�^��ƛ���x�r�sH.Q �yujP�뉚�pX�^�C�evX�ϴQf'�P4�˯)�;G(s���YL=�=���O~�C8�$��7bCc�ns5(֗������WP��1j��m�V�e�g5�M[���!}!��:���ɳ�%Cye���v.���N��#��_E�f��܏9��aP7�D8���h��;Gw�D�-�a�F	���d.(Ms���RSZ��73���p�P|�����گ�&
�H���2��^�f߁z\�A&*�{��� ǐ�6�,�K�He��|�G��Y�n뻈��أ�z��	����#uH�&[��d;L:~�ID�)o
��?)-�a����Rx�1�}��?���WK��Um�b����P�?����b����P�˚:�7��i\]"�,����z����a�^��8#�~�vUÊ�RLX���hX��Y�b���0	���RT���N�ԋ�7S:��z���^���< g0��Y���&3-d��Dd��9΅�LV�g��M�+�����*�C��ϑ�?	��{���L��*���/s��I>��m'O63��1]n�r5@�)7� lp�[�� ��Q��J����[]��[DM�ӵaJ� �̕������hNJߤ^���ߒ�N��c�Y�o�:�,����R��,)c���Z}��k��J�gR�cj�ـ�\����9���B�i���hFT�ע�նJu��M������8�4��ѱ�����{/s၀|MX������Q��h�lRe;"Ef��?B1�Xg2��	�'xU�;��z�?�~?I���fs�o'=g��J���i��]�:=1�.�f���}��ύuJi�%j+��g��[v-8����-
�z��hag���K:^�3#�\(��4�*[n_2�S֎�o��P95��oP�(Y�&#��n�BH][��W��n#,����P](�m[�6�0��qm�v��}�3������/�2o���k[3y�y
H�[C_�-�o�ڢ�8��E��T��R��X��r��w`F�cT�]<�I��R�!���n�iB�rU�in�]}��vY/+xj���d�p�Q�����(�mn�O�^b��o�<��Ǻd�b-|F`�����q/ ��#��(�?y��Z�����M����Lߖ�]��F�l� ��ӸVi�25�^���<�����6ʥ/i�r�����b��rU�E�ԟ������Ʊ�I҃Ӄ�5*vib�z5�X�a��Z-����
\Lx�|��hn�[F��b��}�['��>e��L�N�-���Z���]���j�UB������
�NND�l�q�.���}���'��|x����
��?�Q�դ��fG���]͸Q�7����iu�� �wv-J��8d���n�ɖH�����(�M�Q���J�
:���N��;���15�ؒ���h�q+ஒ>��YMH?����o�<��S-��r[xR�DX�=:�@e �g��vB0\Ѭ/ԗ�d�hc'�֣B���_�