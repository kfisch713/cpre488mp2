XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bs7v����P�o�D�X����"_��o�/��[z��}.4!b#k>C��"ά����/��@����C��#���������i*�����gz��� 1X]��Ѕz$���MK��� ���ܺ�b�x�h�l8�Z_�g���L��A��P����ac�Iq 9z/d:�j��/l�0��oξ�+�aZ��PcD#��`
���ѯ�&�����d�ԛJ��ؔ�$���Ԝ� �H
[@�1{-^_��I@E�W������2�ԀèɬJV3�P�=b��%Yo7#���@�۠S�'�q�\�C��K��L5SV�ƶ"�#�(�O �A�^��Qߑ�B˜�Uyq��-%G�.�"���V�P��@�=�Q��	˴��Y�X�f>Z�&=���|��W���)/ѻ�C�
/��O����l�z��7韕&*_t��@?ܩx֩xb��P^X�:o�h��O��xx���3���Y���G*���<E��((�������7n` �+�dX�%Ŏ+Al �2k DY� �£4=4J�6?~F����0~���-C%�p�J}#į�קS�������8��>�l�#��V�/n�ۜ���b��2���XF9�������6�Q���V�h���~��p�r?}�T~���rܛl��4}|� %Z���� �.t�T+#�-��Y��5���K��A�W�>�茟G=H�����U����@oG_�p��ǨH�lH ���p����ƛe��o�@�r���
z�V�E�5�XlxVHYEB    9fc7    1fd0Y^�Jd}>sp�C(�.'`5��#�3X�oƘ���u&�*������Eƕ��od�Q���� foelS���c�nK�րb���J���-Dv�Q6Ђ�gѵ}��!A|����.p}�i�M�t�FVJ����;���U�@y����;�z��M�� 5tV	��4J$���Ef���Mu��uQ�L](��ӷX�pXY�pd�,;c��>�\Q��?]-���Y�d�lR?�@z_:Y#n�w+��?��>d�^��jĉ�_�ӿ�&&��E��������#� MZ�<�*�M��k���A���J���ٶ'KU��.��V�z���U��ߐ��Y�~��t�7���]mm�����m8p�fM�Q��^�W�L�1���b�'Vq�yw�a���f�aiz�L['������:��PU���Ev���Q��PX�2��~Sd��N�D�i��r�����H!ؿ%�:��F&>��u��-��|FQ�w{sC�<��r��}��ũ.��i��1�N�ӑp�3�!e��kq�.@��~VQ��l�[JMNõ�D���F�����[c�+xc纟��9��A#{������z�T�I=�4�5�e��?h�2L�ȫd��^P��W�X�O�6Љn�/�������"[��pYH+i���R����e�5����kș��溸H!��p��m�I��~�I!ǡ���� �v}C~;��@����c)��"�Y,qk��Gf�jw��V��@�"�����X��즛�=��63H�`)Ƴ��T���D�D6��������^��v���α�A�g��v�5&�7�!�Lwߡ��+����C��\��h^�!���XH����#��vE��@���Z�R�� ��y�d7�cA%N�y�[yE(��a��S	2�:Q�~����ʧq鎁�@¿`2U�A��L��<&E�7	)s�$-��u����ATـ뗟UP��A������Dm��@��'��Q�W�����쏼��żh����3]�4��ʜ�d^ICZڕ-�������=ū�#��S�Kp���_3��k2M~5ߴ��P]_�AJ튢����8���?#G�م�UI�#tk�/������v��>\F���@��cF�T��>�����_��I�ޅ��;FlH�\�e�q�0G�2��nf�ߺ\`D4v�%l�m��,�,5�r��dA�Ov�����;^թ�$�f���'~2� Y�Q�t�=19��O�ݍ��p�?�͇<@�/Dި[�m`��*�v+�t���,���̠��/�@�$��:J��D�D
W`�!a�h膶�����[��O��nr���0���ix 6��%@�߷�̎�/�xM�V��N:
}�A�A�%�B��� ~�%1Y�dfe��+���|ժ����T�[T���]jIA�݆��k߄;Ȭ8�P�'3~�m�����K��
!n���.�eolFZ��HB��<������B��dD��G���Rb���!�1J2p�*v��D��[�E ���nV��w�	ѡӕ25�mD�&�d�qZ��3秽}�l0b	%D{r���J��� m.�*}�t���D9K���W	 P��h(
�彽�����!��m}M�`��Y�{ �V�7*��ڼ��0/v� ��_:��^Je�@�΢Ǭ�[7a�ץ�AIԲ��,�ͻ��Rg:���r�&N����E��;���M��jq3�3�ZT,*�s)_~�w�᥵6P�|�
Z��w�{��PIF��ُ3#�T,�E�O��P��{J�^k�L!��Ys�R�e�Ăw�%���,Q��EF��_�T­1� �V4a�#OqPD���^��@�S=���tx�����jm�[F�/*�1r��+��%�s������;���d"a�S��	��Gd�����Ӡ!1ɐ�*�ѝ�r(�3��j��Skn�x�Z+��0"�v
��r$-{�-׶��(���jWS�iN��p�v!<�7 �ڻt���V��g��SHjyC��S���y�S��k�Db�?��b��{ :�F��1����8�ϋ�Du'aL(gx&:G�PP
�0�����{|���,:�!�o�����N�flsd���$ p0L@���a�_$�YQ�\����Ʊ��/8<E�\od>\�M��QP�O�T(7"����^q��Bٷ�FV�\h�:���k��WYt�f$���1��}���V��mѠ�6�S��1�_鯐Kz<�$eV����Ʈh�����s� h���ғ�*�I��q;O�@�o1�6�����gn����i����*M�lL���-��4`SiLy��\U!r;{0Xj�7�NY��<�A��{`W�o�*m�n��~s�N��� ���}c �}����#$@�ZB>אP]<��&4Do������!��&J�P���Aݙ��g���~bgNt��1�������=v
f�ѥߚeӃe��.��+/{y�MR�g�;���/*����*�I�O
&�ց
drc;�8��7�����P挼�3��fC�!�=D~�?�V����������<$��J����)�qr���E$��m5�^�ޚH�p�����Ob�ߝ8�O�Q))� ���5��9����ɾX����_���Zf(���qӊ�l��#�D�Z��=C�^�� +�k��3�d|Lp3�B��?����w!������}�H"����?�FD��mo�u�]T���2tjT&�7�v��>��4�0���r�`n	�<�.�����r%�Ov�M����A#���	ON�L�ҥ��wb��3�Y-H�t$8�i���W���Dߪ1-A� ��S�O�;�1������^zq�Ĕඈ?8�0y�\�-Eq�V�������WN[4PrJ#`)�P���A�3W�\)q��D�3<<�Z���3�BPZG,����-|�g��Y��BJ��>����9�>�:ʃ����NA�U��g ��\��	Y%���	{��И>F���4Ԇ| �S�%��j;� �e�Gۏ7���P��YȻ�Ⱥ=]-�2����Ԇ�xb5��V��O.�jp�����g������mA�7�^�
Z��ۡK�[$ֺyr;�.�
v8)�M�;(��U*� ���dP]�Y,����M�9���5A뎩���H9x� .���
���͵x=!�����iv�����JI��֙)E�w_c$�� �"�8�?b-N|h�kt9�,����<^���� ���f�Ms+G���w�f�J~������2�{>l�1���ǌ��u㪑�z	{�5����O�S(x�@3��x��4���,p���~f�RLU�J�*��3�'��W��W�$G֊��g�t碗��2�>��� ��D�8����$?:8y6ywmL+a�g���u�nM�O+񗼝_&�[��"*-�%�H�Q��Ȩ_�]�i,�ao��aR��*�r��	q���CU�0�c$�euz|��J�G�-�<�hr�ŵ˚&��I���\�^������IR�q�r�K;�����I���������4�|?5kJ��P�.vw[{a��&�kk��RUӾS<���j�'f'	e`s�Y(��{IG ӓ*Jb�_�X`�&��ŠW�r����2=��9y!o\��}8���@x�p�^#��@���d�j�93�+0nj?GE<�Ў1.�?��Żb����O´�QYK,��a���Nm9�iPۮ��\��7]�Q30���=�T��G�PK��R�����0�UE�9�g��A¨j�j���3�=��c��81��+�?3��X`H_	�u�V�����a�����Ba���=�q�!^¯���b�yz)7u䙻��kp����v��jT0�T9u���F�"�!��:�0�rD�؇���8H��v�����0M��3���3-L� 7��ǂ�r��R��/�D&X��DFq��,[Ab�+W���`�#�ȩ���7�:��g���RN�ޛX�e`6���C2�|f�b�zq��׭_�r��~�E�ø�V��H�Olot,��P�C����zA�ݗ"C����-�N�WM��l�߄R�i`�4���@Q�����_�hIGV���ZI')2������˲�-ݤj-�1�5�LEbһ�1��0��o�'�c�c�PޣV�J��	 �z~�Bi>պ�٭ ��ת>�o���ߜ�J�ca[�/�3����t�3�w.,H���V �P�ÏA�C����鱁��Z{�}��dڕh�Ms�D���3�f�ްB4ɜ@X�������	m����P"��RJ3���䠿��/B�V<�U��&��VX��T��H\=������a����)��R2����+�Y͈��]��V�Y�],�w��{��X�����d	3����k2��D�z��RI��f|�	���3�	�.��YN�����<s�E�m	�y��}�>#��3y�P�ۑ4k��$�)u0��њw^<��S�;i�<<�ї�E�$��ڴ�9Ǜ��"ܕi�gJb'/cK]4�*���lʍ�{���g"8��tcj����Z�  鷤u�T�� }ߚ۸%g�*����Cnңm	��e��"����Y�8��!�~T������9LU��"����e�I@�߷���ٺ�����HN9|�D� ΊȮ��C8=�\��"��c�ş�P��i7����ì�](����B�쎟"^,e���֘��`��!��R���ϵV�z���o
L1cN$G���(r�tB��P�3�l"���Y[T^S����P�?�3N���ba�����\Z���%�8b��iҊ��T}F�	*�e���ҺPk\F�s�{�m}/kᨧ������mpYOI�DZ.W�8�U�ޕ�g�@��B�/��
*�:bm��8��a��,����kK��;:z�n�ԗ��WԵ�0=��m[.ñ�d��ԕ&Aվ�O���0�+P*�j���V�#iW�W�^���*�1	� ��)6=f$�����4\�� �I���$@*L�W��Cϐ�ŇLCdt=���{�s����A�0QP��PUV �����V�������`�+U��F茚f���������ۤ]��ZK�j7z`�a�!��TYo#-��K�>�մ�[8q�Ռ����%;ަb�5��'xR�uH���б�fs'�ۛ��|D�>y� P[��"7�\L��W��G�QE��3=�oq���MMKw�h��.�,�n�
4ч�N����e��Q  ���[���w�v��(}j\�׌�� ��Sߧ`���W���QF��b�w�S[3�\s(�r|�G}�5��������IЩ���j��(+�9Ɩ�+IR�Mr�[�e}�u=?��ә�=�K��Rg��o%�Yǎ,z�Nk5q�ۖ'��'Pt�)V�<M�f�v��-U:����Z�p�Mn��xuHK���õ�^э�5Tl�@����P���YCm8	�e�K����ǧ�;AE[4H ��d���x|�FR4Pz��%WR�_$��|F����]�Ār��t�ؗ�A���~}e�T4q:J d�g�����*/&ζ�Ԟk{�����d{뼪t�2���\݌�o*B^ n���H�TM�4H��Jm��P1�m5dveG�T
s[��{�N���nL�2�U����?stS��kc<8%�Β������Tm�{M��&�����:����}+�^�D,�d�!ܰ��@���mpxK[�ڎo۴=����8��[V%����==m�1yי�NѵptT�(�d���n�TCE�\������N���I��È)I�޲�!3��p���sm)S��ʬ�p�\�WC�^M���3�#�p4ֿ=@��G���<�z���T#BɃ�8�f�ի:���N�&��Z�N��$��`����O��tTN�)տ�%��55� (��w7@'����5{k9�ϴ�*7^��3~�B��[�P; ���ӽ�X�
�/ި�R�2����#�7-�<�o"��gΊdVP� nw����h��A���WNz��������MR� �gopi ���bgfZS�SzB@���A��y �rQ1�;'�%H��e:��o�
����K����Y��mb����[S��K��jd��階\E��:Ж���;l�8G���b�i�O6m|-Br'��6�KPE����J��"Rb��kޒ�2P�P�P�*{J��W��?3�F��k�[�#0����j��J�MV�͜(vi��`A��R��?����wOG�Z�4�^�r��J��iK0]�����[=��S:�>��i���?�K��<��n��В5�D�)�v�x�ӚF;�L),ϳ;�T����&��</7�����r͏"g��㺙:FD�$Nb��5�S[\wG�W���S�m�{Ěe�f�:�{�����,��R���j��d�աe��-�vw���H.MjUxa��6�3����j���A|�}&��v�G��ۀ06�i��o�s�l(M����u��vS۩+���-�w m����	h��f���ܳ4a�=��c׾��� ����Y�`�N-�"O~�{�:���(tZ?m�G5'�|*������>�O�+��b�m���J'�ݗ#/,�����ظ^3JH����Hb��ln�j�ef<�l"�#k��doe�/t|���'����qz��^Q�Sy���Lr�V��������ɔV�}0�vk w̎�j`�?;-�^���,�S����?(�-E��f�d ����wk�q�hH1#qy�?ƪ�V��D4��Q��'���b��y�����L� G�����z~��,���R�"� �>��m?�l�CErv���a���5����ΰe�S8k���n��"�Tt�g'-ԇB�
�f�v�K,����7R�,2 S^W���a{���_<A�a*�2&_��ܖ�����#������6�h_C�-N�vKս-�����
�*���6��v�6��bN�$f���������.J�6�zG���m�@1�ڷ�)W��p�b�:A�k*�c&�"�K,B��,$�lGC�'�)1��Ee��!W��8�	-�3�.�n���`<U���ƙA�h����,���s�4��ci�"�$5�~w��T�ZY�i� ��Ug ݙ��[׎f ���X)r�Pvet*�����f��%TૃJ�v"0�V[h��f���o�ڬ��Ϟ�Ӯًw��)������*����:�r�KFk p�6�a�k��!O����eЃf�Z�"B�� ����5�
>�;m���5�z����5:�qE�f�@-�0�l�p�?" � �Q�V:�'�N=������/�$�I���Q�<B�0��ajU%SW�t��;��A�oz�P�g+��xN���4����S
6qJ��h��Ͻ���g�οH�2������NN�:(�va�Ո���Ax�'�;�}��_��cq�|E���w(�By���ʯwظr��������n�Y���*&{�h�����l�ʍR8	'yR��e���y���g�IyC��W��d�vf?$�uب��Y	�c� �������G��^Q3i?p���v�k�i���N���H����*���SM^�i�_�ր�'���-Rxg�j� �Xs�"�;���iJ�Tp�Ȇ�^Sb\�Pi��I�@	�|�����O��8����oC����nv����e
3�(��K�Z@�J?j|{'����=zC�R��~n�Ю�5��g%�׍G�Wtm��@`��V�T��ο\�4�gR%�Jy�(�'�:�΋�ﵗn!/��r��[��z�?�ۧ���ވ�g`��ؓ����e]� ��k��R��
���f_���1���4��8�w�n���a�������`qt��e �w�21c�$r���FTd�]�(���'j)Hۓ�K�_��!�xB�3���~�`0QyH����d�@��z'TL.�:� 	��3[��k��"��v��o��ǍFm�������o�[5�F�IAq�!�u]��
*~��;��a�9v�����t�BC��i