XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��zlI�����[�����t������g ��Oy�59����%�`��t��G�w���44�A����C|��w=�$�Ƈ�.	��9�"�(U]�CY��$'�z+��C����_��w�p�=s��.�݂ih8s��>��F�����Z�p���	�։V �Q��%.�{щrO��|m6M��+�S�3f�T�񷻖+���+-I���_�����V��	m��+eF�f�h��SDE��y$����A��i�%��K�ⴡ�P��+���}��D�lK$��Ih�E��ҳ���2���N�ո{��%ځ�C܏E�O�5�7Ppt��%���L������׮ܫ̹��$J����P�+��L��� ��M���(��L���&�on�^�k:Q4���R]��r�R�.��F��@L�Sr��fd�e�0����N�Xg��q��،|ЩԀS�w@���N�A����4ixH��ˠ�9�U 
7:�9���m/�4��HMk]�G�w-�G]L���!�������{��:�N���F6�Q��Glv�@��(���%�@��(��8\PjMg[�A���WYz���y$@6C��
Zu����y��ð9#�����OA���ɐ�c.�6z߅h5M��W�#��@��м��;V���Vq��C�4��ۋ@ �$�$�
�D���x�|?��))3��T[�<$�\ܢ�뮵�/�{n�u�ִ�����g�?tcay.$%8'G9���,E�`�m��&XlxVHYEB    1959     920����?̐��W/��i��!���<?���șL�R-�/�|�qU��wHic>�f�M�2��~Ub�Y����]J�,
h�i��7]�oj��e�)�/i��#���Wcmf�a��],
��'T��>�����^
?%/��u�6'z� ����N��Y���WN��B���!�V��&K$HE�Cx&����r��M��>>�#�^�T߆�v��ɬn���R,��?��m���� ��+k�4�\.��r��N�~���P�
������Nkb�����5	��֘)��@ӧ25�p�اL�XG�HG���-�h�������[�]b����^D�s׮�� E[�s绱a�D�]�( 4;���������Hl������e|��#E�S����3y�g֡��)���_�UK ;wn��Xv2D����O����"��ܡ1�o���I��2?�U-�YdTH{����%x�eYa9q�D5�s�ά����a83�3&�{E�����T�#���ހ	E���if���yO�C�m�0����q �گ"�������6�ғY-Q�+�GM騎�=WWؾ�8��֜c�	6��Q��ٱ�����8gt�MEO�����C-T�`�I��4�"��a��@�oҎ��)�0<�(�[����N�4��_s����$Zq0"��ܗ�Z�nh3��C`�xH��&���|�Å��)�U��%��G�)W.!q�Q^�E�H�`5QT]6�cM�>��}f���ڪ|EB�+�b'�LC	��8ARksÀ��+���ר٢h��eԉ��L;7C����:���4��k�v���&�;�*R�5U��q����}��Dl�@s����ش[��[O-'wq��:ȗ���.�Lְ�׿W�b��k��N�ev\���kڎ�C ���T�i�i�(���
��ˋ���u1�%ԤZ������ @E�ͫ���S�Y����K*�/�69�����e�x������9>�`���|)�ݝg�]'o�	9�<��mS���0�hI��fϭɢ2k�QK�H |�-ڡ���Ȯ�.�#�]���bi���kE��ɣ4��-��@_/NWYU�KO������/��n�סO?��QϹ%s0Պ��������@r���b���=pPw��6�P�X��c?�P�[���)v�G'��:�AB҃<��Sh�����Eٵt�>π��h�?��#���� ��/rZ!�?�s_�3�7��X�HN1�z���R��5��6]:>��5�~-kS�]�w��R������<�M |g��x?�7�fsAncU���9O�T�=B4!�R���a���h	p�N+q�ʴ��9bv��e���"�N-�U�\f/�m�YR�ێ�[�yoEoUv5w=I�5�T >�goEdN]jlP��ϕP����L(Tz��u��*�o�n'!<P/���
��q�,��!B����e� VC�z�I�[��.��؝f�&��������)s�󲐢����M��̌LИv��VE�J�����5���V��K���%��@s��v�H�ʤ��G�0XHwݥ�!z��WH�&�v��AQ����>��Q2ڀ�jc]��lž�������@�F�<���:��T��W�����u�)f�E���P���6��OFAx-h��j?����Dv�>AJ�����.U�_�1d��k�w��`u�A)���C��\с���Ț�	'@\���Ӷ�������cnrϏ�b��/�����M�~����#��jޤ�D#����6F��g.�A@��@�2so'4!�#�.�'�S&C|'U7f	�3��������c��9�5M4*�L-���lηfd�>�F	_��t��m���-~�&�{ՙ%Q��ZD�8��&�+F�T�'j=��YT����>���������s�4�����+�a�� +(y	�����ln7&W��Ɲ�N�P�hg(��u����/����"G�(Gb�n�G?�"�V�4���-Qk���6^$�\v�c�h�1�kۿ�e(�#u�V��m�KME����/��x�����zbtB��/<�?}�����5�Q�N���eQ2ə`S�]�貢VX�-����4��Kl����g:	���/DXX��NQ���p�&�n>��Y�*�Ʈ��]\��0O��Á�`�5������ +n�u
�]���#��.�1;��wic3���2�D�����s�b�^��>Ý0\��.EѾ�J���<���xGg�G�u�-ٱh7�j,갟mJ�z@�~�vd$�