XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B�r�O�X���<�՝�=ѱ�
��4;���	b�Z� x^Z�tu�ں�b��*���A7?6~�s�,��qZ�\��m�E!]�*�_��r�6���&905��ʟKa����V����g�ȝY� ��Lz�ě������_��Ƚ�W��`ĂVM�E�x��y�#��%3*���
*��[��?R����6]zU���G"�ő �)�L�e��ɼ��j�z���%7����*���Fū�ݘ <�9x�<�}E=��1Or���WL@ax�~#���u_m=�,��a>7%���9�����
�A�11��4m������m���	�4��C>ď4+�1�7�9c���N-��+r���6��n�&�5}�7D|Z����ld�=��W	�?�3�*~��/�~~L�Fp.��d��8�^�*QM�n}�ڡ�@�%_����	��Te����X��,�����@�=+!�����
E��^�~���5;�D�5s��Nc6b���87�\���P���N-�5��v����V	�X�{�� ��W��+�F]�14J�-��R�<C�B����@��yTh��`��m�%="��3Sx�F'��6���+I��&d,��Nd�U�j�������c�����7)����g���^Y$6�����k��H�ܲ��]�	hm�{�a-IA�VeMwmc~�W�3�~˲O�g&x��,���.��	k��q�c��-!��:������/	yE>Z��XlxVHYEB    3d43    10303��m�np_�`W)S�U��{�I9x�Em�:ZȾW~"3u�t�e1��N�5)��)�l�5+;�5D3��^��M�]ح�p���1�J��p댉�!��K|��o���	٘�̖��3�RB̹�I��ߕ��.��Y�ߥ���H�[O���ׂN�C��/��h
�� |PL���%�z{��?��y��~\�C���}6���B�c���F�V���d�����/b��-s�:�uvi�_�KK��¼KK�W��$�C P��̜��>�U{�$�_�E)��:��s^ݧ���f�"o��^���� yS_Ak_Au-;G�QZT�&=n?�8H�Ye7�[wR.���d��/��G�ę����L�L��Z�BD��.��X�0�"0�����h0�����t�a��������d����t)����Ó�Lz����ώ����({@��V-3��z�1J�]��)�f���d�;1 @΄��~�Ja��gy�I��5s(�j��\�� !�Y4nς�D�AC �+�z�c"*��J6J�tqэK�u؎��]��f���=̏�������nǇ�ϡ��s�r�
5��g�e#�����L��`S)���0b�sZ���q�\���{z,�oV7��n�I�NG�`�.�����M����WR�ᣝX����u\��>�2���*�x5 ���l7#���?��vleَ2������R�,J�?E�^�H���'U�����1��8�^t��3���T�h���Z�:z��X$X�p�~�Mo=��z"���^����Lj���r���h�T^���k�7'�$q0�����@M1��(�L��vX�O֮�7�z��S�n���'[d�y����($�
<��\"�e���'=q����G�gg;h�4�y��"B���*:Z�/�h�F�گr.�{'x˾��JdJ�5�����N��l�?s��UC;Ea�X���V�'䌸	���� ��д+����xS�sY���J#�1���t��P|(t`&��	�Z�y��C䊃ࡂ�'���fas�N��n�^3a��ڮ��{�E]�'�N��t�J���QY�!±]a��H��[�zic�N��������׉
��Ю3t"cϥ�Rd�&�>��0��?+^�K.~�-w}���l�`nH��T՟c�� "��H�>v\��=��� <�V�ʠ?q�g
�S�R�����0#T���w�
�BP�e��_[2�S�_ڰ:�$�e��J�L��;���7Cv�M�`��~uƊT�ng��	�/ ���	�����&��-��2�S��[ j�`ZJ�g�6@��e)_�����8�'��wn��]$�T	I�Nqs�.�+g0�h%�Z#q��}b�W|g�@�w� '�'�F;�v3�th��*�s�*�U="��j<{{-��zc�6��4+5�1����\�1�,���N����M�2�_#F��TD!?͞�G!|�S����T񆑔c�!�Ğ�x)��hW����J�c�;�KiX+)z��Zry�];I��!7�Sk�4���]��M�9��Q�_�{���?�y�|p7I/-���r!M�4��&1xa����'������A�Ų��}aT�N���#4FC��N�>'�=t'�=�8[��:`��4n~�����|��E���S>2�lĴ���I��g�\�{��-��X#�kp���k-�ٸ]�\cKv��|M�[�s7�����+Z)���ct+�;C�3�3�����9�.�@�OO7M��꼚P�j���	�p��+�p�����ƙR^%u�=��2TZ��Ne���~��5�DF����I-�{/�3��,��润�_�i*�Z�<�6ac�)~���X3~:N��G<&@&��I��1:c����-`��ѣ�E�d�Ď�T�Ѡc4M�;�r��+~��z������Y(~T�D'P��]Y��yO�g1��ؠѪ�Á�o����y|W��"n�%H�=�����Tw9%␰�%�;���pՆxҟ�b��d���v[��A���XHC0�P�[���3��t�A���\��Bo�i��w	G�=<����4�[��]t;�k�yNz�I�#;��?����Kz"(]���g���e�O�0���3�4a\�3c��P��g���g���e�/ �m���g���8�#��Ӊ����-���G���yu�,�2o�=* 3TEwuάS��|�Ө��0V*T�%|��j�XbS+�p��|?-6V�TLWDؕ�(��t2K"����1��V�h��A�B{'��y��:0/gK/<nq������i�dm����4u��Nz�ĝ��IL�t�ܴ�����}��ʯ�mt�y�sP2��PQ��ʒ$�L&��(�g+ray�8�p��c� n%�����{�/��P�>ύ��)%p_��(�&/����a�>؍�w�j�$s��90�yfIۛ"��y�ƶ��9�A��Os��|X�	$��(�ÓY�ĶXJU�
��SE7���:S�3ic� 0;���N{��Ư�p�"e�kn:�VQ�n�I�����қڟ	dߓZN=0l9�����^��]F(=gr�&�z�������7g}f's}�%��������/!2!`�
�_{�8W�upO�����g+�W@=*�sxEM5�.�Oƺ��T�H~V�`�^����}O7_���.�4�a��8�q�>h��d,q%�p6��-��8a~5�h��*b���uH|v�br��+g@q�u(�g����TE���,�S����k���K�!�33�D�3�Jo�Y��H���@�'��H�)= ˿,e?�4�x�:N�����_��c������<]��!~6����s���$x�����r��RR��>�|�]��f�Ԁ,-��" �Y<6��l��vS�wͣ���S�;��_�����Z�r"`C�6��<ra"��L��
S�/J<$�{�KC���1��}���:��h�sA��W$��k��7�Y�P�Ae�9=�,k.���K-�M�+�]��Jې�1gy�wK|!V�E��Y�,0�(V��n�螵��cƬW������?^���+��eg�g��y��������)�7�ro'}/3���fnhd�]�ۣ��&��['�H��(�s�����&)w�SgJq�
���>i��X�9�RMv�Zb��v���	2Z�q��)7^��N	夗�>�߀���2��T�r9E6H�S ޙj�^�F�)�ߝ�ѐ!�Wu}&��Ӿ8`]�0��/�V�L���3��'���tb_z����f]���=@vf�G/����4����r۴�"X�J�r���?HH��Ph���xd��6�x_W,R�E�v�3[4�t>7��&y�
ۍ���
��&,�����;���c��5�@������ �2j��]�P�ml���/�؃���^���*��0���b��b 0��K�Zc��$��7�+0��4�wr�C݁rX�8�:�L���R]$���a�y���. :��Ȱ��6��~��rMx]��0�c+O�ô'y#_��r2_K��u����ѨҶ�K�y��\j"�"�p����;)p�Xye���v�Z��q�d;���brue���A{��]�~	���ݰ.�rY@0��޼�p˿;-�q����$�yo���?`���| z� 4XG^�j:�&y��Fw�:[O�^�a����B6�G���aA����B������f�-�%����Қ��K�����xB�J|�5����0���ܹ+��ts�˰�%?w����!?15G�w�� ��y�6)����0e`ǹ���l'��Y>�\2���MAU���=��`�	bզg�f(������� �S�v�����1aO�}I�Uu�˙�6=����F-1�a܃��N��g3
�}�c=�CՂ�T�����8�r�zW�*#�9"�̓��N���J�`)H���Tl,��G.g&&�T"�K��5�q��P�O;%�������/ ( �
wk<�)j���8+0��w�_i^��N��ROa��R^t�[E_��z�u6��R��=L+;�U�����j5��tIF