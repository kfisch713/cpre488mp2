XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b_��瑦<�loG��(̯��P�����v	Hi�p�Fk5��!]Sf�<��}|B���0��~ŵe�S܍�!&�A����� �9��A���:�$y�Y���FE	=Bt]7�[�񒺤��
4Jw)���(���ÿ<Xt���������K��B��l�uZ���Hr��/@�e/�Qp0Y����6��qi��;�n:�t��8;��3*�tix�{�.�X���X���x�B@�4�wx��hx���:���a�����+?"����{�W,�
	Z���bSF�Z�D��u���b�Q��?�Z(/��:�#z�m�M��w����|�w�%�%X��a��+]�F�|$��l�1��L�����0)`wBp\���}m�2r�	�:�N}^+9���x�M��o ~q��w[풲QR�Dr���'(m,�m��TV��������RJb{zD�ʺf�G|�<�`�X�_���X��+;�OQ˝�GG%�I��X�.ܽe*�y��h���L�dq<5��Z*Jb��e��bx�$�r��j;����x+vt(w�V���	{�i��
'��v�f�,�ﵫ��7���
m��'�6��� �?�*���������ͦk��B��O�vJqE�[����+���AXt�KV\��LDz��n���D�=,�ʶ"�S�%�Ł��	��: ؛p-���P�WL.�YV�y;R�*����;2|bL~y�'u��7B��8XlxVHYEB    17b2     880"�mtq����ԟ��`����
����y��+��ٍ1�>__ro�����xH�eU����zy	ɭ�����6|�t[%iΐ�-ߎ�]�iJ*����tۄ4�H���,��z����g�F�����mGA���d߽QmV�P� H�eg%"d�ZNh\���J9���G3b�c C~�r�z�)�eoJ�Uz��1�|����8	���{�y��ٕ�VR;d@�]eV��e�Ȍ@)��&�D[��z&.�ґV�'��BV��մ;C���-���X��lC�Ⱦ�&������Tb����繬�����/�
�;v�/�{Ά��)�VU�t��+��-��W<���S�|�0I1 v��)P����zf� �{�z��u��1��|4�jg75�>��R���->
���:���j��'[�q!�-����E����j�Q�H����b�: �k� ���$�Ǒ��<����`��9�]u6ir|�����W��4�}�l�=~z����l�\_��!��$Bئ���-����m�{�n
���=cN�}��46G���(��π�,�
�7��?��;�h���Շ�ĸ"���1�W5u�eKE.�XW8afi/
]$i�+��u:
@\�D#	q_:�U?�bp�;+���n�
����٥��)�G5s䅽&;!0'L5���`�0wR�ۺ��JB	,�G�B9pD����w����N5х�ݏǋ-?!ί�xB
5�#�f':�^�-�Wvh�v�42���F��Han�>{0;����ʎ��w�F���}
����3�>�/����G�;�<�Kf����9��P�߸���U&m-	b�
��ٔ�ڳ�%�沧VD����zIX��눾�����.��J`��1�{N�J���`�4d���9����J@[��$��~�͚a�t�ml~AӦw�'5(��h�h�r�H��g��Z��{�܂�-�Iک����7�8	�$�{bΫ����� (���U���{Xa�k�)�.c�q��4��u嚞�R6>R�FU��$�n�#�;1��7����h�$��,�!���:u��P�OM��������3�qp\%�ξ��o��^����2|�~{	���V�\^8od��gvZGe�~��@�ӳ��CV�%�:���71�b)�ǻ�xG�_N`'�2��Ԉ�~�+�	���c������	�qU6( �Dq���'o���xz���waQ]'!Jڢ�M!_�
�����nd��O=�bP�Uu�d�2���8����$��iM�Mծa�\KoN�x�����ECz�2
N�W�ƶ�$�gL�-8�{�G��E"I��8��4��a�Ƞ�W��e�i�(�č�Қ���_م9"�@W�n���k?���5�r-��SJ�Q���QضһG�k��'M� A�9����cN�B�<ɕaB���66?�a���G���y�!Ql��"�SȠ���'s�� �W'���g�_ryݞ>@Ne��؇,��/{���ݔ��'<ڞ.�^us�t�eO�y���g�HQv#��H�G�H&���hcK����.��Z�+k�*�ա��Q���aɃ.	� ZVf0�Jv��J 	�1�����of�$��h8�.>,(U�	~<�Ve��:u��4���ߚtT�R��_�]\eݦ7ͪ�u��~�nW��j-���8��`�c�1���P4
\/�|g9���L"M���6U�Q�ƞ�UZ��X��mSh!p�uW��y�4�z���Z�����%{#�_~��	>*O�����1Ұ7F	Z�3@�],9�_�$�O�Ƿpe'�Ш����A�:E����ؒ����1���M}���4'�r�m>t�_/~��otd�dW�|�L/���W#�U�W$���w�����(���:આ {�6-�n"��S�y&�^�*;t�A���]��+ף�iР�$���x�uE�A8{�x�N����@�`-�G�%>�Aaz*���G7;I��A�	������g�Jg�O�5E[�Q�k���f3QF����Y%M.P��`Hs��_tv�QV��b�@�E�R{�8��j��b���a"o�"&U��3G�[�����L5*"������w��~��/C4V=O�	��.�j���