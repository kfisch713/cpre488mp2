XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Z2F��1�a$�;ݱ�����5rrzWa�"h$UAe� ��y�EJ�
i�N������Y����>ⅉ�Z.#�Qd�vy�����Dj��0mD=��X�א�,�V��-c3�X����ӎ�ӭ�9>9owh�>����N�qA)���(�^8����5��Z_��mP�2��q��2�<��Ÿv�4��ebK�ѐs�O��܂
[򱼞��Lj�F����ܩ�Pq�� �Kћ�$:z��;��s��J��P<��ᨊ@���
%hh�F�+�*��ZںQ������� ���S)�I�]a��1M_S�A�-v����01�����@4F��w	ၙ��tQ�ȔY7�o�LEf���p3P�@���#���_���hJM6�V�J����!	�R$������)g��OV��!�W�J�J	�(���'Oy�	*�V� |l/d5�)�_���y������Nse}�\��j��B�����i���>�>X�C��@5-����s^�h��� /���t���O"��S��eL	6��������ĹcY�T��a#k�dE�Ҥ���ʚ��ԢM�j�����r��rg�ʒÄDS]�~�Z��%Q|Um%Vc���H�9��ٿ�Y����u:?K���܌�`�����q�U�,{�K!n��q���5���Z��0k+hQ5&wśM�ԞG�عx7Q#���+9cb�!�o(,��j̈́q6�d�(8G�!W� ��I^�4U�y�1�KE(XlxVHYEB    fa00    2040sx�^'�ن��m�0���|zUxNO{ ���R)N����e�/�ɠ����WF�,G�G���4���D��9RW��o_,P�. yyN�����AB7>�o��5]���PT����� %ъ�C#V�]���ӍV��J0ڽ8��[��m(����5�A�bnsh�8�t�1(Q�Ԝ��E�F�����V~��.�߫g*�i���"�иl��v�R)P�����	����X��lv�<-���KkڑNy�m�69���}�Y�,�)B����D�!��Ę�WE�9��`��q���mJ9�yL�yK:�>]�vz�$�+Q��8\��U
쮧�FW`�6-��������a��f�yb��7�)Qz��/�,k�Q�Q���8%/5�[V�l�	䓸d��(�)_0J)��H����x���˲8w�;��B��S�H3f�y��[�*���Z豇���L ���Ǳ
�Pn�΍	Y\��O���aΎZZj-= �?��s^�6mC�%n5.[:�>���xR�DA]DYø,�	<�>��#0;5��}��f־�TCP�0N�|9��ӵ���sUa��5�������X��!NCl":ހ_[9��p��&_՛�!i�A"��9^'�]f���y�_;I�2�,�$G��Rt����4�q���Y9`4*��Q��ɲ���8W�A�ݠ/�HJ�(&=H�c�T�Ԙg��T����UC"��\2Բ��/���i1��4�w�$��a�R��id�Rs���N퉛�dU^|`W�/c�]�x��8�-߁�=@q�m;>;Ԓ1�v4y*]v�������7�S�ە����#�8�����	籿lgYJ.kF?(�5�z�������z>M�8o�+N�摜p��@�f��f_1�Q�va�P�N���%s��oS��R� �n ��5X�����x�"�p�,,���Ջ��v�3��v�3,(u5CIOEr�Z��jE1A�҉>���=zd,�m#5ٯ=;����R�1(Z����%�q��ay�.�ɡ*:�]R��g�"s5ھ��)L��zY~PM/��7��^�8��̻�6=?��\c
C���+¦��I�Я)��/�V��p�&�%z��~��zM1�b��gb�i�W�\��	 �~/�biK�4�i�����Vyƙ�>N�r-a�2�ǹ�.�]��@6��Rw�,{̶���ǝ-��8����]B?}��hC�_l�>qI�,tĖs��=��Ӄ"H=�؎��z*>�ˁ��_ ���ǂ�̃��ӷn�I���"lDc����!�`-�-���� ��RkZ� ��O�*���"��g����L�O�G���dK���=��z0�����z?�T����_�!��,a�ϡ߉��#$�9��vB�y@���ʓΤg��f�n�n�	�k�)�Z..<����8���ǂU�}Z-Ŋq�>�i�95�$���X��7`����=mu �%���K3��p-rg-R����Qޣ*��_���m�:V����6,4|6Ѫ�{d=ov�:i�6-#h:�がp^�����[����$�-�>���Ӽ�\jc �����NH#}�d�B�-d2ҔR`K\5W��,�LQ	�#A�y��X"�[���2-G��c�au!{$7�xUc*����2m���aLmҭgc�l�T�.O/�͜M�9���m��"DA�f����c 7,�J�Z�p凁1�\p�J��i[���D�}���4Y+8#� 24,���)z�����>O~��HW��ٍ�y��s��8�� �+�Չ`��pՀ3=�.�C.`�-�З���C~��x \L��С	�*+�OWe#�4�%ưb�Ax�:�JHN��=GJҡ
u��%�Y���;��:ޘ�l�`��2��r�Ķ'�nā���"���H���j�Oi�Ut�m���V���U� @��e5 �s!�.c��z�{�����tw��8@�;ꛥ[(�E	|-$	���L>?ϸ5r5�(�$�]��q��慰�J��+2����̾���Zޑ���mJ��c��c�q�������ρ2���ii~Kj������T�q5�+�-�]=��-����c�>��.$��}�1qX8�U���4�R&G�`�'I&\�_�]�� +-6i��~�`����; �.��н�c�b�F]�"�����-4Y�A��m'#���_Q ��<�����x��7Y���m�-�gb2�*���Sg�1�j� >+�;o��#w͚n����	�Y#�u��t>�h���#i
��t�:F]����7g3R$:s׶�-cA����o��L�� �fq#D��8L,��V1O ]��Z�����O�BI������X)m`����!a*�M��x�P������X:\4�K����}�L+�t �Oi�<v�f~��;|����b���I�{���8�[[�uF���N�����+<B��S�;Pa*w��l�U�M��%7��S>�73+~���*��C��Z8`�6��9��pմ5O��T��*�ퟣO\�+BT�k尴
^W?!���d}ٓ2עe#*!��	KV�I�׊F��J�m�.^Q[����sd����D;���MD:���@��s+x�����{ ���*S���a:�uQ�F���d�����i[^>mO(��1j�k9�	��:�B��v
�^>�ċ=^S�֥�s����s�BO���=w���1���a���^�c�ͶA��@�ЏSF��MD�R	�x��Dg��/t�\q���X0Ĩh�MMPS��9�ut� ��������jm�}�wMl�zv��z���S>��yɁd�Ȭ�O�'�ڎ[ه_��Y=���&vL� ����S�N�ED�Gvc�Aim�]�H̙-Ձ�W~65Uh�gسn�(��,41�IJ��>�n�"%cf8�M�2�ј�����ԜTS�����w���/?�l����p�6�6���bPO'�3��kw����swtt��3����!��A
�:E
��]����H	i|<H�(���a��>&<���i�ŉ�lM�B���+R��mt����ԅש�Z�6u�c}+����q~b�t�`.]����<���d�ab��9��so��&��`�����lz��Tnj"���"f���-�\@8D�!�K�ۣ4*v�v2k�)pa�Cۦ�T׫�����Hf�İ��u����k��I������i8�u� ^P��ïT��h���Ͽ�*�k�q�$�l�\8�`Վt\�0~���7)�ݔ�dK���=�pJ�|����)�q*��,�"sZ-����1c�?a?�qd��3��4�+�3��J��8�& C�������*�>�&?!����Ű{��&/2}��F¾w�������۷|j��#�jh�u?<ak9�E�,_:ZS�{���6J�� _P�m��g�p�M�9�E]BqhD�J(�!V�qX����f�`y�f����}���ń��ȋ'lc��gg�c��j�Kr��z&��	��>Н/ݝ@�p��VL�c�:���LK����s�y�ڧ�>� oq�r���;�-�wT���w�����@�/�� � ��`�)<�5l����dl���W�H!D�O�.̢�e�ts��޵��r�6�#����н%`oH��^3
�t�_�w|���G�:�nΩ?#���}����^��}a'�=��i$`��6{*c�x��-.!]q���O���ܐ�t�~"� w�������3 q*@,%%)n\M�Ǔ��I���p+�dʽ�E�O�mlxTg�t���.� �`�X�t���,(U��k!@��5�J�� 8���a+�����}�h_�2	��)x�������@�20إ�(�yD�6�9}��d��:��ii��d8����6~v�Q}w�W >��;�&ԁ���&&5|Դ�G�4̄{
� S���{1��*�3�օ}xޕ���B�`�`r���3;}����t� E�Z�Ȗ�w��ˌ��L���z\Җ9 wɬ�(�yc/�m�;�(!-����
�<f�aRN��
A��˳&WfF�S��[�X��� E��'=�m�6�a�b�{{��Ι��5�
�b3##5)F��FX	8������x����al�߅��#j���-���L�ܔ����[�S���t���E�AϠ��o���O��˷"5�Y�L��"��0n� js�'�|ҫZ���A���E55�t���!�ֱA�`��3�'�ɜ�DGC��Z�.;�LѴ����*��\-@�ݲ��Z߭��
<ȕ���4�L��p � \�f�Q)f=l��c��8&���H��8E|�؀��Լ�1a�(w�CL���������9~K犤�����R���Ͱ�=RD��'��D��9n�`�`fi�4#qH�2Y˄SfEO��ߍ�����r�Ŕ#^�Ͻ�^{ه���P652[��yd��-���X�ĝԽ���:���g m	�I��ݶ.5�Yº���bb,�}��A��3濳A4�F{�t��Z/�{�7�ER�x'���I��fsvQlZxD�Q�N����C���1���YeI���ЦJ�0�;�C�`@���2��9稜�V7� z�mx+4lPR�&^֩� җDڛ�|�����Ƙ����[v�GZ��?DG����{yU�T�"���|���:�f������zw��0
?Aqu���k��C���}��c�|�恻���"}ỽd���5�0��o�0�l��g^/A���BCR�T؝*�&/�~-'&I��y�(�5�p-��6!�
����GV�<���fOj�
!:�|�ENh&�TM��q͔	^Q��,hf�S�Ǻk�_����9/�j�s!�2܄jFo#y?�-;��_�pz���	Y�e��.m���莪W��#6�]����P����c"�{;�o���4�Û� �����&��E�g�s_ތ;�yյ���q����	�	j�+���4�Z����X�Ȭ<UGoR��Ӥ/���.S%K�=�=�s��C�	�Y�S��g ��g5۾�^< =��S<ҍÙg`��p��� �]�n��6^ڤd"%Y��x^�k�l�y���4:��o��\�8vK�01��H*IimSb{@�n�����N��G�ù��H��K�ި�@'4D� �����D�p[#dI 4�ni"*�Va����ݥ�z�k �Mifӓ��ED���4/�b��b$uyT��
Rƶj������?�ޕJ��6�(�v����{���ԜB�;�ҁ��4Q�7e%
��Z��#����؜�Q�U-إ��z�"{�ٺ�1��%�=N�BMH��ʣd��E�I2�VA�ރr-�3j(�_'��񼬞 6B��`G嘂��F(G<�)��[�%$m� �ZQ����|�^�d�U�r����Ph��>�����:��@�����Х��m�l�0Wa�;�WZۦ�U�.�{&m������.Y����y<{��9o/�}ӆ����f	�9�j`~HT&�?p��1��R�V��?��y��@P����a:�x$��P� ��٦�x��o'�~�^ꐨ��GE>�xɐ�R���?x[��Bj�zz{H?�!��5)O��y�ږV��K��t�o�A��_�0ɲ��z}�`�џ+�K��(�B�I����o��__��)�4���C�C�6jU_הc=�����	'7���O��Jٿ���/� Ӕ<��$
�Z�����5�������^���m6�?:bC�6$�呌W������h��=�)JS��~�8�ckǱr��-3���jY#��~���W�f2�~�;�ۓ«�"��o��Ρ	�3E.�(#�t����r<B�����\�3�д7XeM� _|�̀X�u��K�XeyU�?�EU��@x��a������Opw�e�Zs�H��)�~��[YB���VՑBL���B���k�umAŜ4�m7S�؞����ظ\����V;ۚa|~�I�¢�p���M�;X2?ݓ���HKxw�p7.��1-��ҟ��j�f�w�6٨��<�� ���
�� �G��0p�~��8��Ny���K\ͷa��q��#"j/��BG�i��:!(���)m���s�=��l"D����׫�"��첢�	���ъ�|�v�v9�r�Vӣ:�� ����J�3��`�$dw˱�3>��`�#׀�tу�R�#��DG ��00��	r��F��YD$u�q�He3ؤ�AZ���F�轥,j5��w��2�;�t��|��^�g<�E��^O�S�oD}x{�9�x'��R#��C�H������*�����l����"�>�k��Ns�d)�A�A�Q�	� >~�o0�?Ej	A��w��Hg�r3�b��ɕM؆,�P �z�(w��@�O�	���	O�j����z�>�|���z"%%b��h��f� Q�VzA�5%�>�ً��
�R�~�=��+Ľ���\*y= �!��N�;�H�
n�ȽZ�V���J	A�� N����'��Ǔt:|]0���Hֵ�4��L	�E�^?���Fku�dA��Pѭq^vw�9Z+Ie�q��Y`60 ��q���8 P�[�W��#F��9�?y߰��y6*\��L�w(�mz��n�v����@��a>��q��������T�����*�o��,�)�,�ǜ�0�6AMSA޽WcG? ?�Ǳcw6MLx])�.l;.EY�����[�������
T�����՞-�n��!�$K�)D�lL|?c�Ry�
��\�od+1�/NMy� ~�؃q�MT���t�����?�����"�'f��o�h�I��3Hic4u�lP�3��]������Uş�������K�\9���vkA1-������\6��-���pSNK���z�ʧ�Y���_�A;A�Q�Ϋ*�d�h.y*9f��ை+KZ�y&�����MWU�=��0bZ^�{�@�A��w�>�>�WW.�G���<�t���u�����/�;#���.0k��9��9���7 �}F�;��o	��N�43/�Ŏ:Ԃ!-�r�=G��?�h�v���1�<Y䤉��#vs}~�R�f,�D~{@�̣�|����^ԫ�04�_8�B�U�m�w�(�I2f���{�U���
s�!�皣B��#���Ll���*}���7�e�]�9Z1%Y*Z��*�@,cd��K�~
��5��P���:d���%x�5ninP��'��E�m,�V�%Me��ۑ��5#�������ڬ���TP����'(;n�	q7�Q(��W���	�-sy��Z\T-e@ѻ��oHV���5+P��$ئs�g��5�g&0�.����a��1��͞uݙ7v "�5٦�T:+�k�c�ȅ�ܶ�h0֫^Cٔ�DM;f'�a2��PE�.��V<J�S zQ1�±��̷�K�I���� ������D�v�ߌ�����$��-C5ԁg�jh8H;OK$����X�RLE����K�(����
��Z�¨��6��7G��^���WM뜯�p�Y�'>�9��A$r��i�b�΁�h�x$?������˵�b��\��;D'|�E���/��Q���mAt��-�F���>]�%������G�kff4��HTx1��.�I��b^����2�!���
K�yI	���{h�%b�|e�䲜�e�~b�&_�m�{����}�_�� 	�
1}C��#^��]�tF�� /Uc#�I����63h�JuZ.^i*�,����~�W�>�0iT��)��'U�±���Jx�!��$��٤ӭ}�Q��PiC�l�:1��^l�|�x�6n�*e�E�TgڻCc�R;e&f�I���;�υ�tl���ƒ̰z�6��{�G^�B	Y[�/F&
��6���<�Ŧy��A=��,-]a��Z���4:�����v6T��n�ő����X8;�hVCj�c"����r�f\�?���2\$���P`M��9|��rQJ�~q�C���%\�3�;�L�������PDѨ�3r��8Q�*ש��@y��C�/��"�ߣT'V�ڭ�M�$6���ln@9ӣ�k%� �]�w���`?��R �5��t�q���XlxVHYEB    4f62     b50�.ޙ�Ø�yu��}RQ��J/w���Ԍx��Nc�)#r��S��E��N[>P(�u�7.m4t�|�q��97s�-�KL���/0s�c���{lqP�Q��јѴ�e�X`��ܮ�H���O���� p��vq9�����lM����	�.���A��y��s�I���2Q��ab�DE!(9��C;�m(Z"�'���=�~t�d�2�N`ǃ�Z�Y�2&�����F#�$���f�9���^	X��Ϫ�k�'&(���,�(�q��*j��<!9�˰�l�I�Ŭ��Ml[�*���ω0��hWzkٱ���c��Dw~�AEU2(��t|c|6x��ɢa1�]�1�k�~�U�E_�Ɨ� ����Z'��0�M�	���.��
���x��9���rF~x��K#�YS �f���!�Ai���ryK/��7��5>j9fqk��\~�fg ��L�i%xLBh��<r�:Uي@Vꊞϫ�s�U@�Jw(�dY��#:J�6d��@-a�p�z�F�#�ű 	��._�Q$f�0�e�S*TI&�8����dN����q�LM��**�����xs�7@�ʼ2�G�~�~8|0|nEu��rYe����U�B����Q�Z�NR���lb~���ɘ����n=�yJ�?�Z�}�@���z񱫦�Y�I�㸶��/-ͩ�F1��j�-;�ޭa�g���w��rn�t �5{:uB���[%��͎�5i,�p�n�a��6u�u�W]�1SA��ԣH�k�o)��2CG��Z��;i�T\�G�r����~Q;܈ ޤqI����9n�o���r�4�8���z����F�3��g�5����%.|�[}%0��\���K����1���K�9�K�����/��	�X[-D��1���[2��9-M�^UV���.��:{!BH�Ij:.|��u��}i��aĺ��Q��٨.��-��@��[zZ�*Jχܶc�_��T�h�C�#)
��5	4E����n��B�D���4�m����>�J��f{Q�*�=q�P�F|��/�@J̐��*Z/GҜ��+����%����1d�<Q:��;�V1P�\��}��u�r�d�w��)K��I�J*H%E�r��O��r"�ð�	Rb��B����g�d��2FEw���~mn�,�G������4�ٷ��L�n/Z�m9��%��D�����z�l~_=�?�����T���%�w/�y� 4��<m4V��|����E�@3�y`� R|t3<��<d_�<���p��u����a��Q����z���F@����7��4[�}J�m�J^6�>�~V��W|-̶��@;�r�����Eab����Ӷ�'�<NS�	o�:y�Z ����=�"�mjp��/�Α�	�R�B�xqD�tN�B�x�_"�M(>�\�R����A@�i�e�'��w�9�f�n>�Ph��)�aFh���d/��0��a ��_t�m��(���=���S]��s"?�G2a�=��Lљ�v��e�=~r�1z�o����?�6N*&�tNr��$O���_���3��0��q>�̐���)�2���"�h��Vn�&�ױYO�砵�}@d«�M��8F��4�fD�mB�U���A��6�5��\�'�!�݋.�f?x+��y,�,.$n�V�w]n�Ã�̻�"�����d�q�A~H`A���=?�5�t�t̎0/���R]ZW��M��-6����Q��G����D�y�'eڔ�P��-U�D���U�1��P����N�K�)i2~TNh*�'7O�ڶ.�Kl�`��jl{9�S�f�GQC�/E�6:Y��PB�·�9
?�@��v:��*N�{ֵ�]�2���w|ho�5V�I�6SĘ�#X�ޒ�@AY
�k#��x�]U�腤o�$�z�ٰ���W���+��cƓ\�΋3��~\�e�rc�r��Lڑ}A�`
��)��mj��	;B׾Z�]�;o��a@r'��b
4�Kؓ�UX�1$}6 ����m�v�0?jİ���+X"�e�9Ğ�_���۶���nBT��^Eq�h�0Π`����p#�Fd#�A��~�#�&s��;�����`��{��S6�S�n�0G����l�s�E����6�f�(W%��F< ; �.�5�^��Q��Zr��4�7+)�Ju�/l(�nSP� {Y�lߜo�4�=�����ڊ��<Q�0�XY�F���K�-�Y�9���P���1?^���jF\�t$�� NU�Q�I���ų���6�p� yW3��C! ��
�p�W2��u����]iߺ7-�2���X����/$��4�u{>qU"�\7��h�aA@C��&�)rw[�����H��?�#���!d�1a$���p̭�Y�%��w�^,��x'���K�˚���U6Gg �r��M��n��n���h��;L�@k`y��H���k	C2�{s���3��,m��3���Ί�B�"<m#�����w�����M��Z��Yv��i����R��d<��?Ѝu<��Ad��muO����'�⤏[ZpE%����.�#��y)#���R�z�M�K�<k�	e�u���G-5ܲ]1��ҩ:	* �fl���?��6C�L��<��Kf�n������0�>�A����9 &*3�0�7h���,U�=�1��Ƕ�L�5x�]é꠮��l���+[��m����D�j	���{t�<;��DzsB��1z�Sw�3��0Hs���ޔ䞱n��>y&r^++3�t�4��?W��ST��+����으����������!�MJd��CN��V����2���i�a�LO�