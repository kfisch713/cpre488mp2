XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���5o���'&���x�(�@F+�V��T��A�1�y��%B(}�=�a&�$5Lh�F�1=���s%��_��	��p�} mi�ZS	�}��:�a\�����n���r�\��tLf�w���{0Z�C����*?g�\<K8�&�X@�
���$L�����Т����p��%��uɽ2/1D~�δ���I'�]���.K?�򼨡2�$���E�Ԍ� �F0PU+u�J�Tսz���٬��:K�4:P�Ҁo��KR�*㼭��0�sC	u��Z�-Ɵ�k�f:����.��'�����38yy����PߟBy%((\���?Է�t���J�ֶ2\B��V5���OT��&R�#���|lu�r�̛�b��0�U%+�v�hk@9�3"���3��r/� uw)�nhp�Z|��O�.�7�K�)���_��ReEBn��}�c��w=��p\���@�΄蛵P<?��cI�c�U�$�P[N�(d������U?>�.z>�n�����gW�݅��ߢb�$�>d��v�ETF2G���md)n�C��M`[{1�$�8�����c���(A���b��;��f������ǒ�������?�#�oU�f�����I�@� E=�z�Sa���n��|�(8�AQ���(��� ?������S.�̝�^��=il��r�=J����'�TI��"/�N6��~eV��������Tu>`r�-Q��7\���;kA�;1{rS
�~�Y��XlxVHYEB    4284    1110Õ���H��ds�f��{�zQ�5Ɋ��|t��5f֎��!A�$�0{YwvWI&^˄�a��q5�ȂL��|��2���t�S��������f�`U UuV%W�4��9��{fi6�Zo՚����ۚ��d�S+��OQ�U��]w2�z�T�A�5\��,O���1�}�eA�i������Q�P�W9^�"C�ꖉ��P'v}R��mW�4�(L+|���u�l�dO�p�|a̪��:�
n��C���Vw/}��G�y��:30���O,M�6���J�f��L3z��?g@%��U���T����L���	ix�Q��B�I�b&� �у4�J�?�� ��v�q܍jýi���}F��9�b˄%���J>�UZ��q���҂�9^�{sGN�H|Q��� B�@�|M/�)�g��G�JL�����cD���1۟c3Ok��T@1?gG�Yϸ�75������㙆�J����q�tȤ��]�����e�3�����d�z8�Us�E������l(�g6ӹO��]���ļ fT\��~�~�R:/��$�+��䀓����uZ��{�B��=���󍗓<��Z���B?u]$7{B�^k�9�<�=�:,�#UXo�����8T����o����g�8�w��_�M�$�,Y�m	V�����,�����ϱu*Ƽ�\Bv�r��-.��&�%�f����w���<W���`ëS�4{L�	*��_<����$��n�&F~,��4==pB�~�Uԗ�r�����Q#�������~~'e��H?��g�;�Y/�ӟ.j���_���7�NC��aT�j����-���/����vk�^����nĻX�_xB�Ϥ�崮�^3NЋ��|�[|�>�����2`�88>k���+��j�HKL�k�N�ʌ;V�N|2�� �iB�+�ezq�#|Q��h�y;h���X?��L����Dט���SK�yC?�+�L�D�.V�kS�7��v<�"���wOYQA�5��*aH:��EPk�Uy���G�u��憊(��x03A�����2,��`�8{���uZ-vL���=$���~���b��W���X_վ��\7c���6�v���SG1��=�ޱ���DW��U����;[Tj�?�5׺�Mel����݇��F�$b���Mg�Yb�=�t����Y�_L�����e��(D�b�A�۶����,fN���'6.|�.%#��a����-��B�[C�zܻ��	Bf���!'Z���]>�ZƱ�?���{���_���ѢHE�qM���CQͱ()�g(|ED���f��!�����,ak�|ƶ/<�=������yqу���؀!��/}Ct�sj�^��d����KB��A�S�G�`���%O`#aNo�&}��R�HVŽo�y�n�~K������ξX��t�B����s�]<~�q�]?�x�5c.՛U�FZV��8g8�~I@�!(a�5;d5��^* �6�Kf�=m�u�@�4�z�i'~?/�*�f�@&��+N����Ɯ���<��zcu�\��mo�Ģ%�an�:��	���ПP��F�0�~%�<v�X�8P��/\Ȥ�^�q�ZV�� ǣ2��ʮ3"����nރm`�P��v�8���vZ�^_���8����]�Ӆ��r�O�|G}�� ��W��(���;�b{�޶k4	1dØ����}��;�A����!�dk"�B;�sΆd{�1��1�@�|��fs	&X�����SE��+ؽ����u�˨�[�&�^<j���q���o{�+�ő�{�s�D�~�B��E�N�(�Hޔ8��C�lP�0��ѥ�UB������ꊘ;��q��U�<����Y�?ಈ�p�g�h���#�j��*���}}pcD�GV&��!>V����XwwQ#����vPἳ���#=SK�	���̑�����/�!��Q%��U�Yn�� �a}
�_ކ/p���Ϙ���K1����3B"Q>�B�_�0���?t�sc�枨"�������P܇�8\���z��rm�r���թ6˱���/��(�� ���tj_��[.z(���o��e���%/��J�)n�ǉH�?2�?�Q�&ڡ'ﲅ�ŕ¶�<.�i|��N��B��\�m��AC�ml{����V6�-�����o����T�ѯl-����m	Sf	���O�V�l�'g�Zx�9��fvr�Og��(���^D����zw��mBc�+Bbϵ�s�����R�`���%�e+��{�Z���f����-L
�3ӣ}T������[~C��`T��Z)1��/�n�������w�7���2�j.��$'�e��\��� ?����X��ꯤ�*z�,J宿�N�]S>�a��B��s����@�������P�;������R��&y�!��@�'��6 �]�:Pႃh��H�R���y�	t�������b�Ť��D���l ���i^�o�+}�;XJ�՟ҵ�YOX��jo6;����ߎ7뺪%����{O���*��͗үk���:O>Ӊ�J���YI9�}nhȞ�O��fN>����#Ϫcy��	Oc���`�G�Ԟ<��LQ�Z�����n�f�s��X.���!=���J���v�I��H����D����D������Ý����Ș֦`���7f���(-�������s�m ��
s��<��CW6&r�'�e��"�3�I�1�;������>ｋ�gQza�lL����[p�Z��?���i˾|���.�m'D �)��@:�q	���ק��V�}2SC���w���ur�[C-�����x�5�ֶ��:^�aO�R�[�b'2`�
6�D�%�b��"��O�W#�A,�3f	J='�d�%�Ĵ�����C��J�����ڢ����鳢8N�=g�D.�h(K�H��85/p}T�Bj�a��?6��1�2��J�	��ϓݠ��n��a��~�(���#�W�������]'���gp�p��&�\^p�&W �i"��x�H&�Reʶ��cHt\-|<�)�y|�����Kl�;�&�c�;gt&WU����`����C
���Ĥ�%��QH�N4�rKC��}x):LãW�"�1�4�z�~<��/�˜��PR!�m0뾅 ��ԜVI�a�H�+��#\� �C�M#�I\]�{��z�7w!�Y�A�h�%�20A�g~ϔ
��k=z��(�9,X���{��i%uH�X6i��{;>d�?���b{ѕ<
(��F�
G��3fV��7Mվq�p���FN3�fx���Kem)��j9=�+��Yt��R�ͅB.�K:2�e���N�g���c���7�����v"p�(�;�űШ��F;��&�W�B��$i��ˊ��D�9�ū�w�Z�ϵ�0@IE���y�q�|W�8�#���;�Tc�
����-�KѺOP(�Wv*��<��f<�w�����-C��^�c��L�������juA-���PЃ��<J��eևN���.L��h4��%����]q^qyϲ$��{����j���#��}�N����z��o�|�hP�=tҜ+�uu��81��pn{��TD綷���I���~��YU�`ķe�t9$�D���Y#r���Kaݰ_�qb���%bJs�$�[�x�	�؋�Q"�]�묬�x,�p�-�����o��������E�8������Q	�1��*�4E�obBU�A"�bO�ۣ�y��e}p��"�u�>�?v���d���9�<:�v��AE%�7���т>���Y�Ѣ�����۳��ϡY�/�0d�kuz��+2N����gͳմ�J�T`��N�}>:�ҷ�b0�i0���:�v�$Ur~�A�H��oQ�N�,�	@q0��F-�:�r��&pW �|��(�$��!^0�͡�j��6�ٳ�Qdej�`FP���U^�0C���<u���R8��N^�fV(B�K+l�v�M�4�&��+��v�^��݀ϣ2��/�Z,��=7��u��̣S��O��XL	�D�QeO�d�y���Z��Fg���`!��0���s�|c��s(����/*Ɯ=��P�	p���=��˷��2�Xa8]#�;/	ԉ�������"q������X'����Cnj������u������N�i.��f<�+o I���,W�v��ʒ`ͣ�y�T�,'�lt|��tʛ%B=���e\�/��}��,<�!�+n&�S�r�x�_r��̴S(p/=x��5_��4�$?�'TJ��;�Y2��g�����e���tQAҮ�Ob���*
�