XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z��|����GDE�g�4�}k�
d���̀���{p���·�:�',[>��A��v�X}�<���-#�K�x�x:H�-�AH��2��o-'S��_��C0���'�^\VU��63��^H�J�u(�:�E�A3��)�3�?6X"ܝ�:j���s.����=���e� �A�&��Wl�M�}>�^�J�df�x�M�g���z�A@��s��Hm�� ��V>7N��tlnd��C#�B���c�v��V��Zk�����%*�'�� ʎI���y�7��ä��L�����pN��I�0s2����J9%��ڲ�����o���X�r��u�aϖ?W��P�?_Τ�� �:-ɇӎ���r�̨2ֿ�T�!q/2w����آ�qp3�u�[p�fks��^���"�-/�� �!s�,<jۣVP�Gz��&���rZ=70S�*��ǒ^���<7�؇a�u
���pcɤ�cw�!�f�>�G�P��:��ԧ����Кc�8?�h���B�T�a	�JJ�~ٴ��5�P��X���f"�$�ؚ��^�:^"��X��QI%O1�9��f���M��� ��E��'P��6X̅���ˠE�j�����'�ˇ�66T�'��"(ئ�X��	 U5��?j�������Xm
iy�ʠ�imi/��H�z��`ܾ'm06����!�o�uG�KI�`�L��l �I������;�9�#hL��{L"~� �Y���ۃY�'tXlxVHYEB    fa00    26e0_�d�BE�kl9FC�A�rV~���"��ќ�ߢ>�Ѹ�	M��. ���!"+_B��ap�I������ǝV��͊m3*ǣ�w6�K)�	,��R��E�:�qcp�#Kv@\
wo�9��=��u[$�����L6lf��(˕b3�/�-%�ͺ��@��Y���9Te�S����r���Wy�{/q[�C<ld�*\��i2TF����+0�gQ����|-#���\ �W�u�! Ha_N|���.t&ߍ��)^IB��ј2V�� %f����tf#�=�G�zyD�t����)�ަ"�L�]=X�V\�1���'j?�X� #^�O�5��c ,/����������T�u�)a��y��D�Ѹo��ᄒL� �Ed����6 i���g���#Ü����:3����H���Cw����LQ²�H��j�-~�9�~���B�ExB��]ݘCt�(�:˥�N�Lun�é������u��8̝dG�Xa%v3����<GE�b����b8�֦�<!�&p��ˁ���Z�ʖ�Y�s��Gך�I�Eਣ���`�q���8����,M�&3s�I�m�M��.�t*���ߜ�ز ��cƎ�՗=4�2�Ow���&�#eЧc��E�/�6Ok�~��rw)8a�^�����
��ضY7�,��]����)���7��1ib���y��*?�wV-�f�t}��&\Y]�Y���xX1���򥺯_��W͆ǷyN�V_�C��R�>�ʝ�n�t�'u�q9z��f�m�s̓H��5t�;ھAY?�L!P�A#�x�ҞR�Q��.�.�Ka��˹����'ա�)0����S�:@�gkE��茽���M&����D����T��nQ�ztג�lW�a:��w�KWI����ҙM3�6V��'���i3?�2��9H��u~f0l�+Aە����Λ�E6P�
^�T/�L��\6�_�+S�&ޫּ?�G���b�>������1d+����E!��:`d��X��+�~İ~z(�E�d.�fo0�Qi�VҎ���Q/(��[��P#V1m�i���ŔF;i5�?c$Y�,��,
��|4q����#��Y���V�.�,����&+�g1�᧛D����J�9�4R	�G�Q#�$l�)Q�������}s�,�ъ���\���tx7	o(�0�p�d���n��*J���YI	�|��E`|mS�xxtʰn>.3r�0� V킏��i#G�oUU����H�q�Wy�✟�4��z*Ň���-���7U�`9h����k���U�W��f�zp7F9K�N ���T#���e�̈ܨ�n���~�Wu'��"�nz�v�n�P)uZ�H�"MK��W����,�MD�ߠf��D���DY��.��������sq�"���0�&�Q��C?�LɅt�r�XR*K�Sl���c�~IwDr�T�[�Q����5�r`~����ݱWcpN��gW�[���}����5������1?91�:QO=~�P�[�Պ�?'������^�Wm���ꭘ��J�Tj�y���d�����hBF���)�$5��3��+��[V����S�ӯ-s0���}���P�S�!T1��3"�)#C���1�~����*����M'���]�ZN	��X��h�9!��)@cth 1�i�+�0��&���3�'I���e�Uv=<&|}�C8��l���3�/���8uXwj�3��`���l�Y%0p%�"#r���E��0���E����p�Rb
�49=��'0N�3�%�+'��{tz�eP=m�jO��	��?�t׋K#s�,�`D�2�%D{i��k�ӚW<���]�%���T$s{2݈�����>��cu� TH���I�A��B��_]X^� {I�ȷE��ˮ���q����5rb>�B=`Kv[驟��P�
D�+�7�* �ׁ��C:t/vʘ�ԆQ���6��1�v8vrڥd�����T;�2{e�AR��ڵ|a�c����J��u��p����Y.�x����O��^��M:�L�1L�$��G=G���yD�:���t���T�s�#�fj坠�7��%��@c��j�g�cA���3wۭ�cR:�G'�,y�Z+g��Gl�.�[MH���X�!H�u��%	vd��_���Lh�B\r{�%J���{'��v�]�8��8��C��XQX7��V��Ol�&�Õ�k�NS,��[>�X�ԴE��W�٩P�!K2�n|�is���#G�_p����B�4�*�!�N������w�Fs�Jݣ��d�##�c{;d'��N���"mք��9N�}ujc6�w_1����fH��I��E���"����&㝰���h�<���]��'�_�����z����oW`�}�h���w	�p�*��pw2�]�GT�&("}nn�2�y��y9��@
D���S;��a�M� �4���̤"�]����7�M�~�ac+��ol&�P��+�� a+��tHR�z�����˶��]�IH�oa����� ����{�ڥm)%0�oK�����ޙ{��e�w!g�`>������-+��V��1H�X���:+4�,�աM�B֓G���)C�F\�Q�,�W�@o8?�<���cC��������}y��G`��v?��v�2��S:����M&$�sD�&ou�O���!srg��<� ~�����p1NV&��:���=B,�P��_<q"�wG�a+�u�B'��.��n��"��GF�We������q��.g�Kw��L��Ö9pY�|:cGED����,6��Ds�	�ڇ����!4��1�sN��j+R��(:Tx�b{~�#�j�ߣ��}�Ϡ����-�L^-yN ?�B!5 z��[�@]�8�"�$�����У2\\f@�����GT B��i*A��O�Q���yf��ŧ���4{m�:#,[� �S�L꫸� �`�/k��fN��<���9l�z����tZ[��(�WFx��I'��^�ธ���3M��㒚�K��ێݶ1��b�{��e�vRX���i��/[񵃹�j� ��.{^_�9x�,<qۧ�F(��|�jz6����f�������6�}-z�_4ƚ(���N�E��|�����a��w~�xV�7����c��#_��I��U�j,�.��!�o~n�O0r��l^dĸ�F�mG��7!��iy��ct����:I��6�D��
�����f�  2���_�܅��pe����kr�e�8By*E�=���G��~!~��M�NV������ �2�`sv�f�Aڹ����C�ȭɚ޲�$�u;�(���M%��@ZZ[ �>���z���)�Y�X7���
_�{�i���w{�#�X�5��b|@o�>�b���f��R�� ��|z׋��	���S����N =ǽ<���='@	~�����Z,�B,�Q�2�cN��oi��G8�'9qv  �>��S����/!Aq�o�,� S�����[~V/�/]�$�b�D�Re���X�u�Km_W��V�q�������ez�;@��G1F6BE��4�H�_�i}V�I3�،�j{'�w[�ֹ5������6�`/<�mhvK�!kӌs����c�Zq�X��8Ar$,��~�m���)��3��f�͸`O���:����C����'u���7�;	#t�yz��c4ǿ˟#W
oC�1�t�E�j��kh��^�����������0��<���b\���t3�#�xI��&��0KVZY���ei1X&��Ҡ
�>���)<"Õ9�>�%��Q��~;�����m �q�[�M�щĎ�q��In%�4�sy��Q2:����ލ�UꮲL�w�R����cɣWr�km����Gn�t�����Jj 0p�P�,�{��?�b;��F���)�]\�w�z~Ya������n9�n�c���2����Qm�k �ۜk��Z�-PZ����d��n.���!�����.`~�^��bq>!����rXQ�!�7�\cV�
���]�Q�t���똥��	��[P���ؼ��������L�t���u.ۙ*_�0w��&��ј׌��@��N%�՛���Ls:m,�%R�z�?�5�/��ѹ�.�
Qc�$��ͷ��%���!^r(��cb]qe-z��q�5�p-D���0|B��.��Y�څ4Tdң���7�dd���O����&UR�PV����2�G��܆A���<��.7�v�dS��z!CMUi�4 M��PU�a��u�st �������u�گ0JFY�zr&��uKj,e'��a�,��+�O��Rڹ$���� Jh�{�?:��T��_�=|�pK[]�XPF��b��M;�b#,Q����q?��̮�*���A<�7 Y{7��'Q�Sc+Sn�\'�� �p���^˄gm�����LIa�h��3�e`�o&�C]�Xie!�����r=Y�]�N�W��Z�l/��{��e&q��V��h�C$]�<�M��������g����rh�j0���T0ul�4w�З!�>r�z1�gA(�?����~_��L
}�ܾj`�b� ���x���.^)c�^8���u?|4��Mw�0��DMv5��[S�t����Q�ڴ����խ�ߔ���]���S|����O�áUJ�'�Z^X�:ӥ��WGT/�wχ�14Ѹ0�5Ԯo�]o.2&!�9��I&����/�����`I����X�9��0L3C���ue����f��u����bj^V�&�E������߹�����P�T�E��H$V�7���"6�_˨�.;p7�^���G޶����2uKj���?f�m[�0���̇VO`�*����)tN��x���1j�����W�'���-y%�(p8����H'�
�!ǚZd�/��
�G(�w�������k+��`ix]v���)SB@â>k�/
� }��W�+\��p���_��������	�$	�PS�H�y�dMr/!<�d's�p�:\��D��,��A��1 ��ǎ��J���I��n$���ʻ�'
?�q�z�ƗW܄�Y�_�>���A{���Nw�A��/(3�s�Q�o/:��u&��7dV��
MvXm�y�SY��y~�ă�.����7�ҏ�	@��������ڢde9����C��l���Ug루LX��ߌ���Cs�F�,G ��N�Hc�VB�Y���FA�ㆈhD'Y���/y��xG��Cm#g�=����W��ȠɺwQ��]m��E���?X��L�UX����Q6g�MOE(�*׶D�c��jpں���k�m�9�@M���<a��n�܁�;Ɛ�Y�����!jc����E?l�d&&H.��8(��M[����s��Bp�/S��8����c���z6���@r�,��[��b�:��:_m���"�d�vz4��Kx��u��"B��"�&u	t`8�n\��.�E��_��>���)�p�<���#���K�?$��k��(�b �I/����2�`�zb�[pL�;es�{��6%��DD�]k�0�?���&��
\�pL<��]d.�@��9d,IM7���5�r!�,�P�y��F̿�ԛa�)eV,�9���S�S�|'��/L�ɬ��QE�.L�L�յ�F��X�oI
sجO�� ��2Z]�}�e�1���mB-�h4�c�+�4���<뮔t�q��O�	5�����6QSN$\�il�}�k[��P��.��2p[GD\�Η��*�Y�����j-��8�F˥Ug�X���فKX��X�K�CV��i����_��)fiHhr(:��u9��;~�:����5����U�?�_���C�U�f=lM���D��+/^�	���Ӳ��NkK�U6vW��x��/$�H d^V�k|x�J�j͂Ga�,�x��I�r=e��=ݻT��uw�8L7L%Q.��MJ�_�Z;�_�}vr9h4&mza�F���u��v�V�x
%Xh���6���[��e]6� _>Z��/����&��'��v�ū���\XO����/Qf���<�i�j��|{t�ߢ��삆)�*���\�g�����E�5���H��B�����&�uNo>�٨����Z̷�f�xFH�ô��	V� D��[�0dKyL?�����+_��2�����V��,����@ ��L ��l���G� [@p�pfG�L�͏����8GGz���S+��4ߝ�8pZo�.h��Ń0��@�s�wк�^�\�erK��!?O�^��f3��S2�q*+L�Q����?�Ov�I��S�s�p���w]�|���s�6��$�L�PƦ�E���s��v婕,�K(����`�	�ٛ�ӥ��V3{�i������	�����B)�:�r@�j��8x��#)�ï�T�A�4u��e���ڼ�}��>픐W�+QD4��(0��Ïc��g'r6U8\'��9��vl��w��I�K�3d��Q��~�r�����I��΄a�K>�t��z�5�_1�����[�4������N���dtO�p�q��]���\A^������s�CC���5�wST�
w��r.6xу�à�N'��L���}/ ���*�r+v4�]�c̨b�V��%�q���
BV8Z*`ps>�u:T��C�-�-�s�8���:�G<~%Z�Q��n�+}�ш9}�Y���nL ]8)u=Ђqj����9���ۮ�1:c'�*v������t���Ȗ"]t���z���2�2�$�;V`�2�i7�K���b��i���/!k;�61d�W)��ҹlc��H���x�4sؾz|"�K6��Ҳ�'Z��������I�h|ɩ׃6]���Y?�ΗC�b<�VY�4)�_;$vw�h�+�֖'�����:i�յ�̎y
$#�q��4/I�W��?�Mh	�������?�{�@�0��Rv�cHvT�./Q��a���R�05:�=��d�E��)�R�/n�.|,�4z��_�"��#��Jh1y���?%06�٩�M@�� �h�pa8 G�`��2>��9��܂��o"�s__����j�#C�Q���]����uV��q6h�w��S�M�L��z�+����T�jY��Q��/;Qg� lЗ�=N �L_��%��셐���A>���w��t�pW�&~�m�ء��ݛIy��'�̞>�Q`�Ƅ̚Rz�.�*��P�!s(�*tI�/ �lI�7���,���g!����0�����}c/�(kPʲ�n���~J�Z��4�D�[O|ɕx�汝i�`��'��|ƔbHӀ����B�;Ϙ��X�m"N��E���F�@��	8�kA�����P7�-��n��L(�Cz�$�]V�\�g�i���:==;�ǄA�iUw��N<1��2���8�6�{J��ߵ�*j���RL�����WgqL[x8���3Csf���>�=����`^��N�n�t� X���XϿ�!O;��e����n�kg��S͊h��Q�x�����2�*Vl�i<�ܒ����2+ꈛ���3�0��k�����)
%\n��[��`*��2͗a�O�?B����pu��;��6t5n'�R����/砯��h���s�� Zћ�~R]}5��z��2�f=�� *�W���1Ky�)��	�i�3sϬ�6�b��SXΌ��������a? �*������5S�y#7.'#�ҔZN@r����#P�D̻C qAɿ�1&7���P��fǧ`��YL���+#�?uq�@cm!����
9;�/���Jc���� �1��ru�I0�l�U%�D�Q�z`-6CX�O���ҝ,��qn'=�#8"O�t{P8�8�^B����	CjX����*ҞR�`2@�g�����f	1�U�x�!�]b/A���ڈ��������C9q��W�.,��In*�B����j��Ѫ�MgO�����b$��LM�ԧ*f��E��n���[>I���%?~"�*Q�_hİn$��%�B"�.�vz�a�>�'���Or�Q��W<"}�b
��0K<YǴ@ ��_#ܹ���$�'n��~�l��	���x�`U\�m:<��"���R�S�������=�%�<�M|�2�.�9 `F�n�|����O`�{�۽����όI�ڊ�ȷ����B�JY5<W���o�����b^"O\#g1��N�d��F��Вe0��q�}���Mfd`�G�����oC��$o�#�怇�����S��.�&���,�H&���x9k����C�bd}؅f�2$�
k�����]�@�\�f�A4e�τɮp�J	@��|�h��]t��n� ��-����.734�|Ӂ�KӾ���Ôx��2��MA�YJ��4~���$#�M�7��*e\�J�%����
� d����N�{���D��^���S�����iHb�@�0+7��P�dُn�����'�s���H����盳��n�`��@�ioy��>v&Z�3����*�׹D�F�d��dҾ�^�K צ��9@�V�t_9T?ۢJg���I��oH�^�D���8�l֋7L ǜ	��?����̲%��/�p��&qxa%�r�a�q��r�sF���mS��K��ptb2�C�/^�73�핹h���@)Ӷ�~�䧦�v�7��T�zB�>c��]~��x��Y�ҏuҿ!��
�=�_�dK}_ͻ��u�\����'�6첡�>����am��oUmj�zz(X����[u^�ĶN_'T��&�{���u5)��K��&Z�1P�s!�N[f��`�Z�t���y�4e��@��8��tl�rHו�Ј��NUC��)��3���B����?o�V��	��OZ�3�@Ni���鞼զ^�� �InZC��e��D�:	�D4�UW�^����� 6s��*�Èm�7�+������G-d�Jlc �n��\��@�t�2�hE:±��G��� W�7��S���4r&ng�ko}���>�����ݗ�ٰ1�7�ph�%�9m��:��u�{?����ǚ�kaK�=���+{�G-h�)U���0�����qj,���<�'8C^x^���(��L_���	MkO�Q�Ȣ�[f��� d�ҳ>��5Xu��k2��m�A��}��5�C���x�9i�m�$�k�)ᅵT�_O�;r{��Q�	PY�L��Q�x1�k4� g�P�k��aAǄC=�(PNY�� /������G�����Lt�]S�6�dU�K����6� �)�KiB-�m(��Mj��a�6�{�2����ԛ��QS��8�j��#��t,0�ڿ>3t2��n!��l��;�J��{�2�����M��2R���`���`��춫�����
�p�-���2�, R-�$��D͕O�b����e�&b�[?#G����w���p�8��òb��ʨA:�U�& �hg3�?/.�VOEp.���C����_#Y:�!�S�[7�Yr��`�! ��T2�	"ăl�V�bW�D��7�O������"�����K�?�:"Pk�q��{w�!��jA"��ۡ_/#��蔭��_L0"d�4����@�����MB���Xv�m(��9)������%)�H��M�����T�x������U��e�5������&`Yr]�6=� j��X��糊�Z�������#���Iv�h�6����o��η)I���H<U���,��<��z�2�g9nR��XlxVHYEB    7d55    1450���/	ah�yE>��=�߭����`Y��3�[�Mm��f�ˇ5��!|.��E�L�V����tO��Å����ؽթ�8�c����c��l�ڽFn��gJ��~[HB��V�wY���_?�|��&"�6�g�ԯ�f$�k-��8!Uc�Bw���<�7h���G~4��@�Y*4]!���z6���|]�[�?j�C�N��
���(�7�vPe6P+ �]���{FC'y�z������*x��1{G�B�� �T嘓��&1�'L�1����|6�E�(s'v ���&��+���P��ݜ�V�|�r�xJ0~�J!�`�I�z�e�n<��w�s8�h�p�r����)��|'�J	S��@&+郃�lv���wR)��D�y���JDd@ӺD�[(�Cj�((� ˤw��Q(�!6��#E��Rء)�~X�t�s�	o�4 �5A�'��4�������i�zI�`�Ľ��ۖ^<�h
�r|�z�w� �t��w��3�i�>Fu��_�([.�x;������f��a>hC�D�|5������Y��&����}��6�טD;.F՚]H+�3���	�Nt���p���K1����Tys%v�]^��b9�p]`,A��~��z�e�v+�]��?@<M5�T���Z��W�e�V���RLv�	�@y��3�u3.l>|���\����=�*���������b��#����$���q��*6�C��rz�H��D��v�bz�6e�@�C�5T����ڪ�{��ƙ�����Pd��Y��'>ںM�Օ��I'k(�_)j�\1Py����"H���Q2�M��Ҏ	刖n(,+�t��P؃І�t�-��T��X�~؍W���p��r� D���ƾ�Q�
u�^<V���q�7_9v�%�J#E�m��K�AT)äM����(��͚-�ꁥr��T�uv�6��⌔�S|��� �D��V�1Ս�O���%���fD�V20�{M�.�gc����Y@���t����t�e���ּ���l����d��r��3�;`2E��|{�e��p_63�^ܹζ}oa�7培��U|��P9����?Xm�I5�1����(x�y{����EI����X���޽4�FW8v�b8�L1w���(�>�ڏ�uj9��a���3���l\44�'xŴ����mUZ�c�z�}� d����&����nd���d]��[d�!c��i�'���,����Rn2=�(-gP�tOc���
�W@��rŋ�� p^���c�m�Q��E�?-=�����}�";���GH4�7`�5���j���h�m+��_�����w�y���]�a�F8�jO��M���]M�7T�tm a��jDW�e��&�hM<��q�ۂ&5�/��b�u���a�bI�[ڡi0np}8��3������{��<�s�EM�� ��Bo]����z�F�\��Q[eu��j����xx����s#pᙌ�USE��t��zA���y;RI�)��
�L�9O��f�vc�az�v�|&�Si���39;|L͡�Er�]��R=�1˷K�a>B�3�2i �=��C˽���Yc��N���iг����?�9Ղ��q��y^��EQ˶AF�2�bD�'g;7�`�i 
W(?[Ð�3f��}�p>C4��U�#�}���Hy���	'<5d�����;���L7�4fAN��Fi����^j�]���;�3�������NG�����d��a&�4Y�0x)߻�P���8gZ���F�L�]��QJ�����m�ejJ_��,�� � ��
���]��(WTȃ��F8��$95zB�1t>�'](lZ�t��(5�( '[�&�����]2 #���'%�`��.̎�f��)}6-X���G���5����f�c~�o�Lp{)e�x�?/x�� >�Q?�#fvC=-��gI�GFt�8m#b���@��x	��� qv�O����g�A�v@�Ⱥ=,��X�e�ဗ��95m%�_}�V���K�|�|	f����ެH ������0P���`��Z�L�򑭤,]��0�$	V��l�j�����l�ze� o��6��x�� $�Z�Js�FQ�^���pN��W��T(lk�Ƣ@\��-�D��~��8v���
;�M�C>��G���|SFE֥� X�p C\*��gW�(]l�2U&��0Y���u�͵�:��_+WL�.e��Ȑ�[-��p�����mU�h��^Ȱ{��@#�gLf����IY%e��}"����"%���W�,8�eQ�^ծ�-��+�}�o�EV 0��DU?+M��[f&�ԋ�6��8J����-І�DT���S-´<8�rAG�}�A�_��֚\�e6<� �Ij�j��iJ�͸�n�E*2�=�7�0���V"�%V����Y@:����׬_�����Ͷ�fZ�QZ��0�J8ל�."�̅�͆��\�=�ӂ�OO�ȥ�Rρ>ή�Yj"��3*��a�����z�/��M�e�E|I��;�v=>�7G(Be�w��<����Ap7����i+�]�d�"��(0���Y�s�,�~2Xۜ@s�ap��|H����w�����U��Q���~f��q���[m0/��i0�AԜ[?.�G�;g� ^fOO�Q���8���!@�.4T�'�l�@�*蘾6�)L�s�|4�'_��
E�'�L��i����6� ���1����M�aov���jdu�CFSO��ؒ�T�ļXl���5&�������:��} ��S���b�A{��;}+	ٓ��Tڭt�h�H���xX0�ZdAW�=��2�3�M����~�����^n��2Nny���z�/k���]�8�?1����&G�m�^�xe��b��X�ަo :b.?���dhg#/���מW�ϡ�GY�|�ϡH�ǎ~H~�Z̠����u�A���KL�ri{�Q�A���w�U�J\���I��"��1����>�K�_�)b�gL�̠�YG�,D�d�뀲v&'rKK@=�ܭ"Ni����;8�����;��6U6�Ut��Ȍ���/�̧���c�\/�~%�o��4f$�Z���
�D��m�IǰAF�d;{���7��ղ�,Nb�iH̋}1���r��� ���DCN�vD��x���(9���5�W�Zf������~>�A��4~��Z�ؐ�X�f�.@�_l��#0)s��X�N����{���5�L����Gx6�� ��[�Q-��66JO$�3�qz���P��Ok?��θ�u�|蚆Ĝ���4���<Ku�=)o����g��=�GP�!r��93����ٖ1����c��
f��q�1�d{���ɂ/��eyI�}����T��.�.+b{O�:����D@��"O��
Fr��x�)����_�b���ܪ��"����&;���p�eAfrmN���uP�������]�������8�be�,����q���/���w�p�Z��f�����'�|� �=�9w犫o%�-X{�l/�L��k���K�������6�aHyp@h�Y]_�l�T������W&��{Xp�N�������`��<z>�$@�PfF ��fκ���S�#�nv� �)U2�)y�ey� ����ViȲ�4���U}x�H�����K��lst�����O��<�DJ
��K�T�^\���	bC�� ��?>T����x�&X���ag��'3�P�;�AM}�U����|@<{+�h��&<�y�]�����!��]~���F)v��� �J��g/ ��K��ڽ�Ux���;1��F�4�S� �K�I�!#�Dy8�s�ˑ�<GL�{�tH�J.�"�!4����u��507i:��C�9�?>��n/Z;G��h�3W
EAb��\����`Szb�D��M�鼎 �B�8�$�&����l��N�CUѺ�u �>�a`Ĩ�,G 0�i�b��?��dX��L�F;�����˗�#&���M���e�Mf㬣���),��@�]d���V	�W
m5�*[�e�?;��G��|��F�*RT0M'��	����W�tY%t� ؆췴��Hsط��U|+0�:>U��(O䊧(�tm�|_j���~��@�U*O�9K{$Ɔz�b�3q܃��n=L�AxeD弩�K�����
=�c>ɲ�lf����&�����'��9���@!�Ru�R�Č]?-�QY	ݚ$��5H����J����C�5�0���+N��τ~<������I��Hξ�3!����FT�+r��M�GK԰gE�����$Fb�F��گ��X�D>����fHK��˵�=���:�j������{�7Ex�-�2
��&򼓇�l�M����Y��������?�n|�ះ�=Zz�H�B!���ds����R�t,�(�����e+Z����Y��#8�S��k��X�P�`�\��V��$�
M`�!�)��sM	$���[��٧��$���s0=������*�2���c~"�h�?�d�[ԝ�2P'}�ۣ�&���h��	��p�_�#XN�n�bz���E����9�i�m#� F�_��(J���B�W�Y�R��q�I`��������c-�{A!7AG� �LP7���#zA���ٛ�F0��e�w�Al�[���ʓ�e��!���c�h�<�\�o�#�;��E�0��Ni|#��r����W��'��1�����=�{9v555ƮS����rS=z��`���f[�	@��IMus�������S�	�ޙK	�{G�x�=iG�2���+�^�ze�/qx���yb��#:/���=�$˔�u�6�D6��uQ~�WA����P	�|n�������]�*��ި�F6?�8���=7�`�?>a�7�Np�=m� ��X�N��l��9Y����X�Ԕ��$\�̜[[Pc��9��$=Օ��O�e�e���V�|&��T#��o��ȿ�ݖN�k�脮una�����|u�C�2��-�!���rHޢ�����	���A������X��,��&����?�­>����V?�1� K,�(Թ7��cS�͇1�i�!D�c��d���