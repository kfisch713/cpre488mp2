XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Cx59!Ң>���X�P�d�5���wJ�^T(2��T�ƵCǅv!a��XU4dx%��kvh��L}���f2l�k����^I
[dCFZ ���kr�'�
:���� N��tgD�^RO��3��kE��4��H�s@���A6�w�<i�P�c�T�x�g���[5>U��fVA�Ҳ�wU	����I�d|�_)A���&x�DuO�A�:�m7nV^˭#��yc�<a��xQ��	��k�ze���]�$�S�ۘ�;i���J�ѕ_@�8t�H�+��2�C�I�]�/v�rl�=8L6��Z���E7����%p���VT:��z}n�x����+\"��H'������K=iS;��r|�Bnt7h�0Ɠ�Hs!��>�$G09�$d�L�6�����پ8vl�a\�m,qU�U��~nb:n�3Ҹ@���a?��,x7s�[q�(�T�@ģ�j�����o@<�J��T�jh�cܧ���FVa�yҞ��b�CYj��^+�3�����qdK.\"�vN���q� h�8<q ���W��Ӱ�8�P)X��1������?���y��K�o�nx�V֙:�^+"}�D�*6e�p{_jb������pS�%ƚ᱐���v�W�����)�pO�*�{k
4�Jt9����O�I���)�Bϻ؋7�$��U��M��/��8z�u5xݝR�	�ܳ �թr�
+3_��m�z�־���>�4�n�;�h5�*��QSG��fQ��y�uӤ�FXlxVHYEB    b087    2540�z�7�x��|��K<�[O���S��Uw>���Cg��Y�qG��Ys�0���ȥ��W��5�ť�;�ݛ�WO�j�"��a�^���m�L�UQb�8e*V�NI'�YA�˿�;c#_�	�Xƶ���{7�cT�c��������*f�h����x�=��:��B�~#�0�MҰ5��ř$�(��kU��Gj��~9Xۮ�78G@F���+=��e @h����So�G̽Qgvhg&C�$���h]�Q�7�9����J}#�%�b3�zpj��,�º&�V1��Qn�#F�\7Ŝ�( uɫR������4��cߦ�({{��|�������C&j23�x���	W��sd|i��za}͎����_T�%�3^�d�3��3?]��=�.� �3.��f���)j�X�bm�w��@Z�=u�SPL	�,"kk�t��̍�/DUs	/%܌���_P����8�>���9>��oG�g��ǲ��;j�I��G?�����~X�A�
h�%�ܭ! Hn}��DL����
%y҉r������R����1�,\
N)��2�a^^-�������e�f�T�)W@�e��Qete �f �@o��._
8ú(�v?L�(�mR_�R���'kq���hO�����M�Iw���Sf�`\�Hy�
_�O�� ��V�:��lL���#���ٺ��.2<p�c��NJ������F̨!豢���گ����ݞ�p���z�U��k�~l��19ᜈj��/��^ŧf�y̲ܩ����.�=*hN(��aN$����j����gR�F�'�>�F�%R���f[�@U �3:������w"����l���=9'AA\�h5�έ7ӛ��+Y<=��v���Zi���\��dw�䕵&d����>��9^�� ��a�sĎѯ��QLJH�{����OB���y�A0&�����]g�xj544R����*�:������Ca�:�C2&��\w�J&���M�;58��K��e�u75�hL#����:g��]�:B`�B�!�>:蠝0�$ ��;-v|��d�4�<��D/�=�"��G��|����K��Z�ޯ^'��q�E꒧S 5�#ח>�.��.�3b�T�ތ,�3
d��bo�/�%nJ��.�L'9�2�y�>@�=M�-��5i)o��-d�·$<��*[��:��k��-��'�C������}5���\���I!0�)� D�#
O���'��(=�ve ���t�~����߽SIzK�`�?��e,��!�o.���4v�.�8p�B{��[xo���
&����OkF��j�2g��b�_T	JB���Σ����C�O-�� ��]����������V��V%C�
RO��4�B�ZE�΄��C�u��JE!t�?*����M/�u�tⴢt�\�Ӝ#�N����\7��9��~���;��Q���MW�"S��-�d���T��L��w����rߠ�>I,:ק�L�}�	�6t��;y%m����O�k�^Ti����7�!D��M8��9ܬ&?�Ae�e��6�C��Gqh���|����g%��4��~�M?��Jj�?��Uc�\��];\�B�XZ��AL�}Vږ�t_�e���XX"OŨ�� �� �n��ْ�4��~�_T�Bk���Ɖ��KI(�]��YYg�l�ɩ��7Ù�q�۝�nM�&����g�ت��骈o�2Z��ؕ�e$K�S ƚ�t�O�`����b�Q/�6F�O�{]<R��{p[��=�t��3�Vb�愛F�V"{���j��?}Z�P���{�-���2��6&?�{�:�heϳ�;��0|����
��M ��~��	ѓ,{J�䲊�e���'���Qkf�/�|R����ˠ�Sg���"��
��
t�R@�CU�t;�8,(a����2���Ɖ�R�3/������vQG<nMP��Y�oa�W�t��55b&�{%��b���{�'��l��H�9����%���J�FY{ܢ/��JnՂ�M��"�ť� ���(�#ڂ3RvCү�0ڪ6���R؏���q(_�ǂ��!�H��p7KoOs2�3�q.p���=㍚�L��LN���R���ۊ�nW Iu��WT
�	�(�Jv|�P�4�.��(j��U��@�~s�3'��'c�P%�	xQ���
�B��p�8��9A>�ݭ��'�"|l1�>��<�Ov�r(�)Dn�AŪL�oի�*�?�ϟ�Mv�<pp���foO�ؒ /]�}��Y�4K�hhuL�7~�s�C"�G�[R��h�X��tV�pd�Ć���_�2��p9�p/ܓ�;@�C�W':�V@�B�8��$��s�%�����-����/��g)6�.��?=G����Q	�=��b��IcU�����}��,(מ���,�Ke��(a����GH �З��ً�r�t3��<��7��/7�#�e�����>���"K��){���������v{N��smsZaz�J�1�
�Z;(<ⴇw=�d�/X���7�^�(ٌL�CD�Xey�-�
�o˰��fm�>T��^G�iQ*�e�p� uŁ�$ę Yeh��MD�����[N�3F�⋯�z��l�ZW��O��|e��n��,MVɭ�^�K��ݠ��M��ܓs��x�"�S���;8}����G�?k<�b.��BXHپ��T:��*���6ZS6m�t�Y����)p��%Y[�^���XN����}���3�
no8��dc��3$b�D.�E�*�na����+��hb���Ty��ɵ�����OS�'y 6�e��yu��$.̍�"2�Z�� ȹ�@^�Iq恽��	�ᾑ��SY�q�N�I%vx�4�H�lR? �;!\��=�}H�on�#����O��b��Y��a?�P��������}M曙���d3���	�]P>j��D���B- ��4��B]��X��?�&�OXk�q�;��0�Ƹ� i3%ˢ� �̖�P���I��LZ�3�(�i�އ�d�� �Dg5��t�K�X�@T s�F��0��Q��ے���A�C�ވ���U�.N����t/)���Pߑ��6���^I�j�=A��sN��pZ���]�\Ҽ/��=9d�@T�5�]�ޒ�'�uro/��g��W�z�A�J�w�ل>��CYt�ː�2���qCy#����6�"�oR�?�u?0������L���)ܪkzs���l��pjpZs�>�O]���k�T���M�uo���k����~0�S� �A�@VZ~-�-�v�t:D�g�{���,����׳~�7�1���������f'�?�:��bNW"����%~Y�(\t-h���I���g�Iǿ>�W 5DI�"�`h���~�:4*�X� �3���
q��Z��ŝAs��y]Bٿמj;��W��v�t��p�&�ﭒȫ��]��(���coi�Е�?EN���2��Uڗ6vh�S}���{	2BB�Bы�����؄��f�=��c��&L���\,<�̉2�q�z�b�&�0v��]*í,RF5�v����E�OI�	PƩH�����vM@D[�@�H�-|Шgv���n<���FNZ�t��s3� 
�5��|E�S�[cU >��{�^1��T&n��2�B1����ˢ��rqz4HƉL�6
��x{ P�l�����c߹�O��f��Q71~��w]���+&�P��7&͉P�Q���Iҭ�Y_oI��nU5C��[_��a>��� ��Fpb)L��'�<���Nj�/�%pT�9��T�m�|Q7?��g�ۉv�`k/V�8�؉���cdz@�C�dю�l]����:U�C>o�CF-k��/�l�\5 ?]I�ے�y ��@<\�|�Ez�pឋ^�[�>���_ވD�A��$�A��d�"#_�]�"������6��$8ʻ����Ȭ�k�0�C=W��~G9oyj@��>!�����F"[�e4�ў�_P��c�`��k�)j.���R�rgs��37�~����θ,��Ս�:��a��,�w ��߽R1��AH�(C�-��^>ф�B�! ����f��G��P̿?в�Y%j�V���3��Zs&U��)Iv��<�lA!��æ�0ڧ����]N�[�=�Hu�_iȬ�F�mwA����)q��>��n�|@�b{�<ҵW;�l?]qC���)�1�`�6�}��ȑ	FP�5�s�j�}A�q�|-ܡ���O���#ys�Nwh����p����x�wr��� ˴��\V6�<����hK�>������<C�y�
��c��1^K�&�f��^H�}��)�|\��z3��C���"� F��Ȫ�s\�;Z�3b�+�bZrKT�_i��ot�/}�C97q�X��um#���ެ�+��DHS0�m�@h����R88��cU3�2���x\�FV1'��ҟ ?/����m8�!��[o��0*Z�/JA� ~�*u�@�k|�=2�7����1��ӵ��`N1��w�͙ү��Ȋ4w�J�va�9���5�5�! 6Dl��|H�)���_.��jx,R�A��B�j:6r6��r����3��@�aO�AC� dd��J�
нR�h��,Q�������9LV&.e��b��g��S�=\:��C�����籍���N>�"���@�Jg��O&;�߹i@���G1�C��|�b����u��> Y�O��C�I"��D��o���3pA�p�H��q�T���Y]O,v4�{]Ӽ��"�&�ʵo��#D�lb��U��od@��ވ���.� ��q�E����/zQhK�RD� �G͐_U�jFZ�蟩>�n�z��!����Cm������]w�ka���(��f����83���8����[�i�����>���!��g�v�R�H]���I,���U3�x>��(�A�o�W�Q���%��q3�!�8��3�qSqВVH<����8�(�E��8:� �|)n�8��s�mm�4����_G���ƀ�r���Sz���|��vܧ�;}��[?NSC��oКx)0qF�S��x�/9�@˱B�C�|zL�ȥ,����&O�� �U��m�E{�9��АF��,� �~?9����4#�Y0�Ey��<��T�r?@&��4��M&ԏL^)�B3[��xq>Uݳ�јi��F���J�v}�p]�"�5�ЛX��; ��4�����:���B�^�^ �T��/ �4�� 8�/%�^���Յ}lE��/�Q(�릸S�1:ע.cDB4�Y�q��4jl�Fe|N����Y#��QB�6w�b��U"�T����U���u��G�tƱtED����ΡL[��1�s���@���v����$<r@"0@'��pq\�n���R�u��D�|�A7�c��B�2�Ϻ����x�إ;j�{{�*��N��� �R^�ˢ�j�UX�.���C{��Z79�Lrv0�(1����u%��p��bKuӡ�H������mȷ�g���4Q��z�+i���^u�D����c�v����M�},���K�pJ$"O������2;lڢ�ý��ͱ�Iϝ�S��� ��
��R�M�N�?��ݼ!�g��V?��G�"\�,&k��ݏ�"aG�jD^��C�bJӕl� ���T@7�G�.�>���R�btT�(�s��0uP��ё3!Nze3���5�c�,aK?X}\ܝ�%r�1(�+F�u>ŀ���6�xU�T�컼�7�@�U�v,Gv`�*�	�$������,d�z�>�0yK�8���=�#V0�܂���s���4nPm���ph�m�g�����'�s��i'�������ғW�؁:C4V���3��?�4#;_�=JUzz1]eG�a֐��A�����p3��<�ܬ��GqZ��m��W���t(K�K=�l���d��ޥf��(gC������,wi�ӘF�s��TS���I�K�����_˔��:������:C��(d{���i��:\��Kh�Q�#C/�T(U${��R+&��p�8�ߎ�^,�2��\H<���z���~�[�zq��+X���Z��ȼu�8_cWV[1L�?���b�7��{`k�{6�w�qƁ�B��G,!=zl|��Sƽ�/P^�7�Y�!�	ޣ�@��(�L:�?H�f�2*z���S���1󃁞pt�լ��e\)�A�FHM1驖������'�x9�e�,iԋS��
"��Vup	������T����F�Z��zVjl�vPK�9����u��c#Ȕ(H���������2��C�]ǌQ�\o-¨�i�վ�\�`��~�I��0�� ɓ	 ��H�:� �#޾o��y�Δ
�Ƃ��q��nt&t�1Uq���«����P
��}�!�mүʓq4P���c������qfW�94����\����r^^�1�N���*�Mj�����n΍��+�zZ�`}_��]h{�cٯ/!���r	�1��sa����!-�q�{��1s��N	+�p�A�q��I��7���,	̇�2�]} ��OfL=Wp.I/13"
��Dz���U S�m3�0�,;���ړ^��׵����f����m�ϊ�8YAn��	I�Uy��l�WxP1� ��=DG�it��%o*ƔX��h
�>�n��fETʺ�s]b���4R�m��y�!�L����3ߟE0��c�w��^�s�P�W�=E�<�;ٔ�z��tz�w��^��򢞡��o�u��F1���a�>�
�vV�0p��bR������<��4�p�-�itx�7��
	�l�0b�⵻�ں�/�z��r��`C�L����"0ˇ2�WÒ����P�B���>g5�p��?g	9j~��m�I�1(Bzk#Ŋ<u���"UHo��a�;ձ#T�����CJ{��F�O>H���C'�0�����m2�ف��X{������� '���4]#�)޷C�*z�������1NS!H��6튑�X��j�qy�U({� ��B��3O���B�B��tI��#���ĵ�J�O�%r|/�F\~��w�q̡��^��9��>@�-�:u>�hP�� h��Y��.]60隑��� bX\�U�*eJ����Pu4%.����uw�?���i��k
 vp	�@� �qw	v֏���K�v~�=kG~�R�Ì���#[�W��q��bJs&�C	_]kh6�?��uT>C�������4I��1�k�Ƈ@����rZ�I�w�uQ%vB�ﲝ�=��������7����̿�M�O�4�0��c�@jY��#kJ� d*9�{�]�����/92�݀����P�2�'O:x]=�'A,��I˧A�|Ӎ�wG��ZWj08�d�,Ӫ�w&&��?�@�vG�g����AyJ��\1���xvM�pyo�.��]y\��>�.��V�ƭ�����$,߮��~>�/n���`+D�� ̘��,��'�������ȡ�x��9��V�I�Cݳ�h�5��@����+ELH�
_��������ķ,�¶�����x�~A"�����7t��K![t�?g��7���IGS+�������l���^�48�дU�!z���Fl����^�h=����/��~2j�E��ع/丟V������6%b��ē>.&mϒa�`�$�#&�� �zg��Q�w��+q�@i�e�l�Ĉ����a��D�X�oPa�n� �k�I�̒�i�2��R��
��~�W����ִ%�:7��oѮ6[$f�j�
��؁0 ��w��*�˰S��g�4Kl�E��}0���i�A�$UD����W����޽�4��TYvn��	�"�N��Nn}gwF K��#���{>'�O
�Z�[Д��K��׬������A-< ]]3!艉�ׇ�P�&i��q
� �����P��w����92XX7W���qI�c�v�4C�bB:�K��}��wC��>����y�(/,�dv�y�i.K�g_n��2D�z�@��E?��r�V�j�%�����K�a۞=1�ï�D���`Å���oq-�_�ٹ������j�=&��#%�<�T@7�;3��bQ9���=���{�|��;�<KT4�k�>ܹ�}�����a7a�7k�����RQ�P)6�x�S���6����5*����ţ]W,d��u|u�?�<г��fk�o���,u���B?#��������y�ˡ�5AԠ�$v$<*��TU'6!��r������5�րc+h��P��ӕY�F��J�ş� �z��$���F?l��q���8D�jO%�����Dx�jr�u��>b�Li�\� �=�C��8���1���X�a7�LM5�O�Z�{��+� `f��&��c�%@����� g
�~O��w�
Æ���"&��l�/�/�3䞁2 2H����^�MX��7��F�B��H�%��'�krLX��	������E���xl���q����2�v���O���jL�uKɐw�����F��c]B뻎�BJP��yU��V��-�E0�UO�m;*�@+j�dBE{�f�r��sH�d���ݭ�:�W3�,M�H����:qq��c�cFlZ9,���U�� }�(�8�u�t
\����Ʈp>�簂��xA�#"�:u��r��e�dZ=����;�k�Qz�}�5�b�{UA�T�]���z�6ɞ�l�B�(�5��K!>}��'�(p��H�B��X��.�=�mN��e��!�q��rN�����U�\��ziʊet���5�߳!�g��7/Z��˦����L������qGR�[%��,W !-��5V윊���L��$�$Ű:�/sZ��;�r�s�|���X�,��tƹd~7� s�f�G)1|U7B��؞�{:��L.�S������{Ui�5{����HS�:^����.���b��V#V��:(��*ޡ�S�S(�?�����W@5��f�h���	��]K슦�L	x+�W��;M��g�VY6;���"�(j	�<�k��4�ܹs��bD��t�8�+�x4+��h��4�&6D���`�b�\J5Pv7�IM��ff�ǎ%X!��'\aU�Fb�-�"�U�R��࿡9qa�U��|���1��p�xE�[�Qx�/NAYJ��s
*��Ł��\���s�RBƔf�� `�Y��N$c� ��
*vz��ʨh�Z�/�y�#�Z�?�9��ol���B�tGĐ�&���u��(;��	��ɡRh@�3{����c���d6��C[�V���5�&�zҠ�ų`tѓ�E^��*�����u�g]����-56�h�1�Єy����k)e��bMBv���
DZ&U[n44��μ���