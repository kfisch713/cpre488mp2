XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ڏ���oB.�l�(q�@���� k�P�rX"v+-��&/���"<�1�"�&p��Ĝ"�IQ;�	��ti���x��J0��B�G����
�+:xH�@��NH��L��)� -��+�^��ڬH	9"�RB���*T+�OwW�)��=���K����U|
mJ6�>��h`�>c�h'$����b��`�u�߯��pK!`�W�œ����.?V :`��/�<C�����D��/)�z��Xݡ��(���H�(�G$`����Fu����}#*g=�ds/Uh'�U�.�cT�`���5J� �R���A����;�`ʉӨ�qy56P���Υ�\I����*P&��������Iȳ��NpNtUG�.�y�(1}�m@9n�> �p�H�D��A�ou���\���Q꼱=��"���o��KI��|V��@���^�o�x��P�y�k�'VdE�;X>��ၺ�ɕ��=
���w%W�͉p��W�x��0��_P���v�n��p���B6*����}D@��ZGYgʸ�wǢ^x��(�0p���� F�P3������g:�+tsF�M"���F��f���54��Ucjm
/&��t/�uẅ́ɮڞ�W4,%�`�>|��V�rW�Ni�4V�ވ0:�f�}��u&�6��
���B�vn~1TU
��)z���� �H���J�j��b�9�zt�V��F*^�J�ԕ`�^��O(*�3i�&����bߖ��M�������e)�'/I�R�0XlxVHYEB    1853     810���rƿ�� � ����_��`��}I�'g	�J�N;ӻ3�������\1c� oj`l����|�ã�Uc	��&��E�<��Z�)J�"6[�x��~�̌���N\��y����L�� [�J���vתn�c������&�*�Ax �cb=L�J
;����m^�3�9��h`P�Gۼdӽ�����v��$H�`�����7<�7$��������Kt��d��p,��EO���9M/��8��\��Q�j��/`��6��" ܻ�(J��-��d�����y��}����� 6�Ȼ��ПiK ��}�A-�{��������{ڞ�q�)���5�X�G��Ch�T1���_|�:�X��,�n�M�ؒn�&;(L͇�Z����WŃ|RA�1�0��q����S�w���j��sP�p���1s͸林��O@ P��BUe���S�~Uޥ*�mQÕ�,I�n�L�0Vt�=�w�ߌl�Q|V璻/�COmVl4�h���p��PR����k��T͑�UD�I��c��u�yZ�̡�����Q��p�q4>��F��j`a�`"S}	���$P��)�*k ����3�_�0+3%�5ґ�s����MZ'ڸ�������%:��d��RW}u9���F��zg�t�<Nq����A2��nᶶ�R@��W����W�3w~���wD�)N>T0Z��;��p1py�r�aF�:�~a�i��L_˘D��4{phoѕ
���(Q��L�������ǭk]9�Ǒ��`ȉ�;ك��s�h���TزnK����ŀ��*�1���֔23V���쐋��H_�jj�,|�LS	��s3�{��gZ�{� \}�ۿ����ʩBؤS�Z0�{{jQ���J�	R�Z��/V�tc�r�_
\�r2ٲ]V\Z��55{Mn�?�6c�K������Z�IB�%+щ�8����vO˹7�P�� �T(���X$]�냑4��EF����1ڂb�n���O���Q�3�@��P��oA��O.�o�Y��m�=b��c�z5^l���OT�s��<�m��Ӿ�ʝt�z�5kI�����:D�A�> �k\q�`L��O�ܲq�ZQ-Bp�g���-���gr�$��f 8��#�d]��5���� ���M�>�%�zۯ����;��������g��M[�����3�E4�)�!=�]�U������gX���)����S�,��Ngh������̹5�7�\��j(�	�Km��kMĘo�[���U'��7�4��թ1yCiT���s�Z�h���:O|6��<���	���@_@&pK�r��˶������˪�s/��!$������������b
�	#^>�k�����U����	0�]>ʣ� �B�_ki��j��]l�*��@S}@��\�{��P�R2)��B���Y��4O~V|PHiG��w��~:��m���@�t��q�N ���u�D�f3������U��x��6���h������7�LS�"5�R0���|?�]]��������u�c��3�w�,�n�R��� 
�Z�߉5���A���[��T��M�`|�W֊��8�c�J��z�M�3�FNi$3Z8��E��jP2ov��+Ģȁ�^���a��	\�hy.��y@���b�� r���i��ĕL�L<
�N�p�$�M��2V˷��J�����0�귞!�w��/��"ϗv�&T�1B˳��֗������T����k���C�Pz&�)��w~j�4�}�Q(����* F��$<.TK��<�7��߮}���1l�z�١���|] A��V����r�9������@�[�����>��k�,�~����y������y^�PUVB�v�cZ�»Ҿ��� 39���+l�Aw�^�(NE$�����w5�h�.����"� �즶�1��ԇ/Н���K}
���U��#�?ͼn��W�j���H��s�Y�H�Z�����|�F|����