XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����/�չـ�dNuU�9q��y�Y�)�ܐ�ܴ	�6�K����T���a��'�YZ�H��+^;dt��Ո��@]�XA�%�z�Yg$�U���Ku�/dw���N�|Ђ~��#�uD�Y^��\c�%ٺ*�U �� �l3�tP���Z4Mr���\;�|�$y��>��6ߎ�z`7����og�`�^��rD.)���f�{�JASE��D�b^8ݚ�[����ET5ۨ�����ܕ��U�6m���d�)KN#¤�?�\a0�_t�hN�B�����r)��#����7��W��!f�?r�l��RL���D��6�����Q��u FVm��:x�uй��C�v���'Tc��1�/�J������'�p���-�{R�S�4y%� �f��?c�3p4�6��&`q�*��8Ө�e�ѥ�(5~���Y��ɣJN��r��n�:l�Z\��� +hu'?s�Òg�B,�U��At����5y
��\�����ɍ!u`~S�bB��H��i^3�gr�P��*w�:����7�P5���Y%��"MG��"�8c���8��^�	�*���Y�ż+�7�P��V���-������v1�c���p��a�9�T�/r����J��l�3	x���8�j�ˤF�%����}����Ë��Kt�y�.�It�Z �q�\PBc�������#�Y����Ґ?�O l�X�HŞ��� +��ɱy�0�UֶjXlxVHYEB    95d3    18d0L�F�3�f�-�����p�#޼Ii� ��ķ�\W�p�r`��݀,e@@����2���>��#���?#��EN���e���+}�i����<	�{g��j�xɴ�rj�|�u!o�t�E��^^
��?e�,���f���ڜ�s��\�ϔ���;4bfC�0a�9_uD+��BM� ���v$q� �p$����eW)��h�kE��W�@A������q=�4��;!)�W���7��ޟb[��|S�]�_#'_j�p�DB�K��wRu6�J_
��
Wj������Dd�1\:I|�F��@�\��Y�ǅ8e��fk$Īn�2K���$ɆˮVV���QHkv��z��Sݩ��foBA�g��'�8+A1�Vk�d������ڧ�1T���>������["�������(%��׾���n�j�෣r@�wgSA�:�	Wh�J�z�!�=J��Ym�1����}9�c[�ׁ;���Hʼ�f=��b1G�����n�pr�JŗC�55������?��w;�}D��Z\ۧk�����2HӃ0��$���|	jOj��L
�.��U�<�-O98F�,lbeƕq@�Ȱ������O���bAliSi5�
�`vSG�?���8jA?[�:�/��R�
ٍ�!Ty��r}T%���Ҫ��Cةv7�� >F�Lh���uu����^%�?�A~ ��3�z"��A���W06��,��!_���C2���i��l����T�o��ʭP؈��ʣ���5s3��Z&a�r���A5���N)&<���w�x��[�WW72��{��aߔ�/���W~ὖ3K�]�Ҷ�'����al�y~���V" f.�=]h$NX����^־���J�≁����V��A�8G��U�g+ )�LQG9��N�h���8�V��FM-~ѥ<HC���Z���e����E0|nM��s�(�%x¥�O��j
4'w��X:Ve�ᘭ��c
���8_R��� �$ħC�6ZJ�p�A���N���ql��m�6�
K�p��5�9:�tU0���U�XwO��e�sw0�<��G��=�V���o���+ŚWO���cqه<�)UI�\=r���Æb�W\e	����!�+T��sl����� g��	ѼIi��?Ob�P�p�z�����A�� e��+��/0@��T6�!rW8�yGH��3x��T:A&߅��#fu���r9��(���A�����N\z�އ�b�8�7��=�mf�T���RϐBJ�l��O�W��l�y��U�B��&��,8P� D��jR�/>�T���2�vPՁ:E��%V�����A��i����e�(�����1 3�yz�9�-Xf�3�q�9Q�XW��\��IAdU 0.M��4����wf��=���i���!�SL��F��I�j��=A	���K�,��H��i�������"��+`1�ly�%��:$�4��S>\�����Xdk���F��U7#���n��<�z�5��muzI0?��8��l��=}��N�#6�N�Ar��< �_6^�������P�.�C���D��~q�l)�8u�P<V�t��d�2ِT�-u_]0��>f�;��3k�xZ֮����i�豅y_>���
{9*�1����yCA�ǴL���r�4GHzń=�t���?%�dU����o�����dl[;��X ������~���J���[��pL�q#��c;��YSH�W�HA�@{��c����v�2\/�rHd�<�:�Ut�τR +>EO!�����&%�����f)g��:�c��8Ƃ�P�n`o��	�v��:�����,oYk�Mur���`'�K�a1�z]���dm�V�izm��j��K�����,�����7?X=
��G|�e·Ry,���� ������f���.��ģ{��@+� ��hP�x����Y'@W��+y�,���,�fyBi��t���4����������)���� F/�WFb��y2��R�@Sn��<^�b��4˽�i�E������ʉj`�$ej�N���F���ز����x���e/G(�>�N'��{�⭂�
&���&��@T��,�Л���r��ma?�Q��#�������w�p����;�}S<U%հ�à 8�����԰l�1\�M����O���JǶ���,#9/��+T����wf��'�[��%���p���c�a< ���ǈ�S�OE;�a�L�8�	�~�Џȍ����e�r�m�'�K'm�=1dW�}U^gB�y�X9��,�+4K���<u�yfu6�#� ��`55-��Ўss�\o�D�a[�]S{g]��ӿ�N*����5A���S�)Q�H�E�PmFQ-O�.��M�W���T"RF�-[�@O��6�
�� ,l�k *)dnb�w����3��58u+tY��q^��F�������3���v09nϑvbGw㴜iX�W��D�����*��r�����c���ux��m�G��@�a��y���onq��R��Bl�g=�E�VkR+���+1u�\�����LlŎH1�PH,.\����SK�����m���aS���cC�J��d��6Pg]�{����W}�{1:���ŕ��R4���`��9��Kt+#�S�K�ϧnnX����z��x�M���id�9_�ލhvW�^|FK�j���|�y���o͘(�YJuj*�Q39L���q_�����+:�$xO�ansJA��vN�R��2'�O�Z�HA {̀��Ϋ9�eT��o�Б}191p���3Fio���O�E�R:K��?���.O�É�#i-�^�ih����L��Ъ0���h�_]����b���y�6���ʇt�U-?�#�25�zH�hm&q)Yej�[ӫ,y[�"~`y'n����W=��r����r�t�`�t��>.�̂m�⳼�����3+`k���EV�C"Y�<�C`[���1s5ê�u@�����o��C��ea'��5*��s�2�@�(����c���Lw��Ip�ɕ�ۅ��sy�I�Ü�@�`@�B~��F>i�`(�z�mjs`�"���I0����;(�Xk��83���dI�bo{�]Y6�^�wK�m �3K;����Y��������P�����enj�v����#(��L-�imnk
Fd��N�����r�=_���f+ĉ��(�<���g�G���Fen@�B�yX;\�Y2�l�J��$&hJ#�?Y��좆�c�).��E@*�GX`^�$+7�g���s)��(;<� ��&#���I#Ğ�U�^F?�Z&�c��/�a�]4����mcC�3���&E+_�u�!ؔ��fT���.�I����P0�U����� ��6���� ���It�C�L7�(�h�z�0~(�CSr{�3��Ҿ+�D��X���Z7�	�D܄'s����#��CmV�Uv�"�h��	F���@�	pi9���K�"���81'�\C��o�(%��)�Ԛ� �����-�?L������#0��$u/��&V9� �ɬ��|CRr��c���ݼ�r멍������ʾ~�oi��N��F��^�n�0{E�\�I�c-�1��SR�N�����օ�rh,���(�Rźh1��?Ч(�_���)��ܓ�K=K��*�#�y�ֶ�ܤxat*��RC��R����Nʛ	?V\�%~u�����L��'�[^:�ܢ7��Q�yN�DƏE���i��+ܗW่�d�~�xѻ�.�/j��l]����֥IR���8�b息��lx��g�~Codp���qeWt�R��ήd����C��i'�������fW@%Zq͐�O(�i>(V�l�P��M�x/�~�y@ڄZcyL�$�������(k��Teݖ�]Y���CrJ�h��@/�wCט�$61~ӎ�^w*<�^��oJt�{/�j�� d5'�&\?���{��������;Yom�/X�K�ݭ�>�%`���S��r�8�kp!1@mP����5�$a;�rq#*��ɬ�)��]�8�p��:?�M*3���%���.���cB�u�<�mn��u1FC���)D<��������#��3�D�W���
�c��+ I���e�È9lÜ�?��q4�VJxX��9_{*4�����3���A`��ؐ:��^��2w15�D&�����(���8���X����%����k��q_�i�z�����e@��������2���pH�P�Jq~ۥ�j1~�Y��fpok���X��Q�A?4�0�q00�xnK���3�ϒ���B�e= �m5{#�����r����G"����^Ƞ}9�gN/��F�)^�����:D|��$��I�n[2�A$3ӣp���O)H)'=�*�j2ˏf��(<9�lH�(�E i᛬�J�}"a�sY�5־��Uφ�}��O1]�!�jԟ??mW�_Ѵ��z<��<y|]@�p����O%��b�� ���,ێ{�QEM[-�B�.� �HD��!T��EtT��=OǤ�+��F�jB�OI���q؁�k��m�*�[��M�����h�=�a�5r>Zo���dG%{wu���J���1�<+'	� 66�!;�%5��c��6XЧAD�CK"]5������J���Ό�rtA��1"@�b��$�x�V���wQE��R��p��#�J��!�H�kQ�;bH ׭N\��TC-AXc�,˹�Gg��l�>wLV��-�
��_�am��bv��Dў�Ҩ�Kh�L��Z�Iz��'�ۙ��P�;]�{��è�k�&���͐�s�%�k�Q&�����a�GVQ�����zX���{�7߅'��v����x^X��*�?���虲����iנ��w����}ߡq�����{��HxF��PP3�u��=�!M���O�Z�g��f6�X��05:2\�rib��;pRϥ��M((WkJ�{�`V� 4�a��n	K�X
��Qު�O�ui�ݒS�W�`d�РQ��b�M}��$���o҅w~�傡�&_6��ٰ�7Mr��pK��&N.p��5�61j
��G�?�J�۶�e��M�����t��o6�u7�]����w����ǎ܉�IP�̃j�	Ż]���LE�/q���	��S�A� r��ʇ��c3v�[Õ�sH.����,iQwr�e�Y+'n&hU��=_"J�c�'P����v����YT�ˑJ�F�\�A�\�R<�g����;:���*���{��qe�l��@,QtQ#Xpl�p,ۜ�a��ӽs�d�sT�;ʴ{��l)�^���x	p}U�-����hՑ��<-Z�kF�������|Tcc���#S��Cus�E��C�l�^$H���T��ߪ\�"�3��s9�4�{�5�!��*����n�ìvuN��)EE,~<�L����v �s7���[� i�9��!=��Mw�<��������,�mR��;jŠ�L�W�ij=�wq����a����L.�fۤ���03�*`�7�"�qu�6J��N��;#٫��0��x�ٰ fV��������i�=��p��̔�����6ս)�9<P^s��0�^���_�"*p!���]�a�N��5���&t����C2қB�O��ki�ǅ�+2T��l��Q*�ba:�����t�|p�����d��o�u� ��!��BlM���3Fŕ�	��vQM��蟬�p�s��B�{B'��U��7:�H��n)�{~�_G-�R�N^+Oڒ�?��2*��#�w58��836����D]%�ML@h:U����s8n�Lh��Z���yO�'cm 	��Ĺ5�(f�g��h���fq���gê��z:��kt�2i	<�x�����%�5�e��"|侖8e�d;�_p'������-�?3h�We�dt4���<)tS�V`6��
/+	�X	�}�����(��o���w�{�|>����D�Ȣ�vQ����ת\^lMeX#�4>�XO����Q#�PY~ը��E	���-ޏ4ݹ\!RWI���tٯ�)�\�
Br��Q���l�^uV�`9 k�^.�}ǡ�I���� 	�A���p�=�sE	��9�������h�ET�f"C���&0���C��V2�$�����)y9~<}]��%
ӧBY������s_=�U���� Iخ���Ow�tE\��O3��6^���G3���ȴ���E�;�p�Q3^/��,�!h�'��^��AҎ#'��r��oj�@+Q�u�ؑ��