XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����&Y��a�:+p\��q���x9z���q���(�<I���IRA�RM(濍Ќ9'Yk�T�y��0(ƚ��ecAV1R����z�tk7������BS%u^���#�Zu��ߣ'`I�� 1�ƅ�݇D�`2������y'\�VB;�a�|�����߱*��$�خ ���ur�R<ނ��˪�N)��1�i�ZŜ�V5�o#��RI�bbRT�T���%Mz�&:%�U�܏���u��z&�s���;�7w~�^u0�_�/QY廉�f��;���A�|zM�y�6��$�MY������������Mho����X�&7�c���䩀� ܊���B	�66�L�}��Q&���l��� ,��n���~�gℎ����X��]q�ߩ�� 	�(���fa?���m�?��v�cC��F,D���S����}��g���L�vA?�ǝy|���g�Y�?M����P/!\��MR^b���ʌ���N��/�dD�xª�g�P����%��n0ˎ��O���/��������W�8%���k~8��"6�q_қńހU8�R%õXek���Y{C"h� ��}�!F�������i*'��d�'HF�^|�nXZ��O�-�ە�G>wL�=�0T����GM��^��Z1�y5�� 3>Z�&D\=��-��X�8P6T�?�,��s���Z+_/�k
Cޙ.�t���L�3�����z����,��υ�-��Do��`q�૝����#B��XlxVHYEB    3a46    1050�Z�,�� �O��>w���o9�y0�*)�j���ϓ��3��-���SZ�N�IL���Qj�x��m�����39�����.�Ƹ�|(R���f�wl͆��� ��岾�pY�H���%�4�	��O������uZiB�����0��i���v].�*��((�_b�������l��fl�E�O��O����J��!Y����{U��̕���»q�̍��ʘ�a�|�s�Uk��b��1c7�;��e� ^um���ѪRi5{Dѫ��c���_I�_ꑦ+�X� ��u����Y�6���҉K�7e�s-�mm����>�p����BZ�����vI�~�ū���f��>m���,I��9-�t;N��x��uc1�}U��X!��p�8xݼ�do�0a���jkl�TґC����*�=6r62�v ����g�(������wK�k��%�k͜�>��F崶5-w\^���*ĕ��]	���=6*-�� ���>�5��_!�#�^
Y�bQ'���L�5҄~{��}P#�M�|#|�U�^ ��j	�=��דi�"e�
䟊K�̋�n���飣��7 9a3v�5�+Ah�^���;�%xD��M�9I6�K�=6.<\U=������qF�y:Glѵ\
�eH]+���~޲Wk�*\��o�$m���a|`��($�-�k���;�Z�4��;Ė��?t)���	�~�8�lM7��S�$��Hו�^l2�?�	����� j�/��?�f��U�Wc��	��M�a�~�Ϝ:k�a<��dWr\��ż@�q�'�?�*�����X����n���RۨB$a�!I
�l:�{g8�n�'�T0s-w=�xOY�/2��Pq"eb���F�H�񜁫��-T��`��gyd|eQlT�^>�vB#�J��X��8
�����a2�%L����m�ɭhbQ���D:ˢ<f�g�|K���^��.a�p���e���#FB#�������2����O���ije����p�()ޛ���N���MU�l{{jNl[Z1ĿB���*|S�R�ohHeCX+2	 ؀�ڢz�/��^	��>`��-G8�1��mb�=�|�H�/��	r��..d�NZ�̫��i>�5�Ս���:�؀I)�"oxm��"�5ȟ�UuZ��n���X��[�����2�L\D�%I"v�T�߃���X6Ž�Cp[E?��G�jH�C���ҏ��S@@����di�����V $I0��ԝE$K_|�K)]���1�訌 ���(ͩ�P ��6�n*<pVVZ{t��)���x��9ٱ��=)ś�;�t�L{�������@ �}���$��߳ f�ݡ�F�[��!+�>�mc�~S�	O|�i�_=5S����2�dO?֮I�Y&�n���n��I��Q�/1$w/�9�3nTc��Z-j�j���V˸����ŵ�?�?V-��t��`ƭ�|������ڞ���Uy�I~����;����Q�z/=�i�VvKۦ���]H�*���}�|s�Ȧl�;��z'��8��x;���ʴ�|ּ��ru�C�b��}�8t� ��UT�iMp[�%�DH=�d�y���;8b���GPg�ŏ'�B�:#��O���Q��r�
F�,���ɝ
B� �*.ꎘ<Q���ւX���h����u\͘���C:��>�S�Rl�ar�U���I������9d��~���t�M7����J��5�@�m��A�>� ����
��tH������@�EB�1w�-�nJ�ijC�aR�4c��p�����p��w�y�2����f{��SNY܂!�p T�I�O�xԲ(G��'������ƹD%{ᛚ.p�(IP\�����r~�S7�^�4�2���ef������+���J��W�m�ȝlRS��S����Ȥ>����幜�#�i�`b/�q��M^�U�̀4����ȍ�ZQ�so�����-��£�	vI���Qu�����u���K�=Iph�)t�v�٨�M��'�G'���I�Z{��u����7�	��P�J=o�=fvPnƋ��y������;�p�z�&��,YFg�JW4��iU*v)���\��LQO%u��S���j�"�s�{ �ڟ<�@/�+�t��$�]�����@���Å�i4A��C�0\"������0���� �8��H���Nx�
��c�|��PqPh{(儑J�E�;�o���^�f2�%�h�����b���$F�:� �yf@�:�s�HƐ���=�[�܈W������g��@���/=�>"��Vw���;�����D
pIS����=׉3X�F	�t�)��!x�O��(y����QZ �L@
^�m%WS�1�:�i�y�=(N Sfyc��7_��_C-�KТ��U�p��Q�Kj�^K�E^��p��5c���3�0^�'�8��7p�-m�k��j��a�:�̱�<e���7m~|k��zs�VϠ��g�r���v�H�䎯��q��%[Y+��6�)\��5�G�ٹ��l�l�l���\�Hk�m�(;΋�5sJ�vmɨ܈���y4��X���2z/�8j�􂍝?�H%[D��i��G����G�Eg%xA�g��,}�$�Z�)�h�����|�{�r��nD6*/����= �VEG�������Ї�����!�hH�FРz �4@���`�x��/��/債�Ȕ�i�H�p��vℝ�=zW,��}�-�<C���w��=[ڍ��)�p�vI5������&#f�hN��e�=����@[�� S�gC9��.d;��-���-s���ؓ<�J7?�}���_`Ң��p�nڄ50%Yy�M�'�z��d/=֋r��Hc�",i��9c�e�5�R{�jc�(���H�7`Ŋp��
&S�%6M��+&�r	[�b��XVk��W���Ge��7p��]*?\)�������� �*���1���d��+�
m(��6]���ΦK���H���Q�Y�p��������'X���G�=��<[��۠R�=�j��'dq�>��y�@$�¤yx�����������7 I=�/*�x��DKt�DVl�;�E��<2�R"F�fSjQ�����NO����Q��)��3ԵDI*ۈ��qW	s(JuU���d�ޏ����!���+0f�~M�~����`!*&ͭ)o��k�:�ƫ��\(�"|(�=��Vp����{����/��
g�O���bsa�8�b��w�1q>)z���i�/ܱ8������1s�5G��rz譂��[C��h�\Ř�6���5Ղ.t8hs8P��$�:������@ ��=ej����=^��iб��PX$�;��i�?E��O��d��5p��o�Lqx����Y�~�hc!��6�P�"�L�p�T�_c�9�����U�V�*�Ň�E���nT�C�C~��zC�!eB�|��x�a���6:�0Z!�"p��,�c3����Ej�W��Ǹ�r�c�������� vL���p��&�R��Tn}�ݼ�׌^RZ�$Ξb/��3ӈ�"O�f�� ��?���4"�;[*���ɒ��O�L���k�9����'SES/��=i�v�4k	��Q�({�;T?]}\Э��F@Cr"�_U�p%��/�(��$�(�v�Z�xT3�*�>k��^/:��������&ڐ�5�l���#�'9���#��{cRkJS-��!Y�ޖ�ƽ���O���tXR�����Yع��w^_n
��nS����{�$5����Ɖ�l�aA��lLwt#�L�6wP�7��.F��Y���A���X�0�	m��ǽ,`<�Qnb�PT\L"1��^
�):}"ﰸ��!�P���T���d��*�8Y�Z7t����t���;�W��yz=1X���@� j��:����xby%�}8�]�i)���Y,�)��1p�V��k��\a���<-?!�,Q�zF�9-.�x���ff4�35�O�`B�V��ۇ,���`�+dV!�*[ܔ��&�|͓c�h�4�Փ����3��}������EI.���<����h
���]�żN������Q�k`�[j|