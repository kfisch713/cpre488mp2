XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������Yb����N��4�A-g�α���I�����~���6���*=K��~��1yF�_��]�v��S�Y�4�W�[B��v�x0�� �m՝��5���A����*k*^H^�If{	�`�^ub����{�kd����}@F�W��3W��:-襘�=�Np�i�G��U\o	��#�a�*�3ʺ�:t���1p7,���on��>͔D��e��ϴ�{$&��l�T��d�=m\���R�n��hu��1�f�U8��3n�t��"ۖ��,K,,m���}�@P���c����]�T�¾��c�ԞZB/B;O߿^<E�R	�_߅�TR��9d��a>��!�g>��c�W�Rl�W����O��M�f�5I}�{X�4���L��!A�>�ĂH`,L���� ��9@dQ��x�-��@5����c���tpE�*>��-]����C�������P^��v��E~t������M+8zI�	�����oW4���g��ǯ�-Z���R�ѹu�7�uN0�	8�k�_������VkC��d#�~7�`���[b��Y�+[.��L�d�K�ߖ��T�:�Qh(�>s�$�A��5c�d8���㚹G�e�h���s�rf�p�?�nOD����X��������wc8���r��UϘ$��Ʃ.sT׻��AK�ʴ���pnϬ�@���r�����n\J�="-{� ��������P��J#H���J��'8�&���� ��x�(F�6K9g!0|C�XlxVHYEB    fa00    2a40�ct�3;�xӡ���и5r�I� ���B��X¢"Ï�"<P�ohz����(W?�+=4br�H���w�a��ۇl�5��'g�<��1� ��,a�׳���<�3����QD�tKB�q$����N��\��u�m���Q?�ے�P��W���j�*v��5����S�����p�F����+�1���-�b��F�8~�J[rS�I��\d�).�RЗ��	p�mnmHM��ThS�d�j��n�#�N����|���)�P��CQ0�b"�Ԑ��-ҹg�Ij��o ��uJč?Lh��mx>y�OŮ�ɂC�US��ˢn��}����!AWm8PU�x���i���Av�hl�	�:��iT����P.�����.qh�����M�]�
}>����%T`B��p֧7�E)5ez>�".d�A�	����L�x��]Y}���S�x�d�<h�TH].�$b���4��V��N��V��)����-�� g~�2R޾��1��c�T_Kgz���&Ρ �+�&����L�Ud�K��{�M>Eb��A�Ml����� U%S��5��,3���
v�X-14�12hr�^!y����WmŻ�e^��o�r���M����H\��O�����.��;Eo����ƻm-̖���o����鞟�/�Gw���Ϭ&W�Pf�b�/b��D�e�7�gm+r3��:T�uL��Y�
���*� fsŦH�Y�q4-8�؛Be����c��e�?�R�jm�Z)�^`9��ַ�Ps��t0HԦ78�y7�}�Uw��.83E�����8|_F�z�[��2��g�u�>SCRT9 ��!��]\��p��6���|V9&
�L6!,���ӷ�1�|��Hr����;�k!�D�br��W�w�"�[��a�KN��/p2��p��M|�x�Cp��+����+�,�pb��P#o����1��8Ig�����}k�$�q.����a�M��r�W;P`���yY�)R��V�_q��01ɨI�������\$֍�%�p3�����^�����5�p��Z�&�]�(�U5���Ƙ������i����	��<��]��������;�w+�}�?��/T�t��!Y�4��e��s��g�D�� #���{��#92�d���"��g���p<���ր��8ݠ��w����O�j�4Wǵ���H�W�Ì��r�Ot�,�ڙ*Z�P�4���5�	��1_'�P	����{i�h_�E�8�Ǣ%��G�I��U���j�P��p�*_k�k���;i��
?E�w�����m&B��zL�"�~��%~(�v3����5C�2���V��lu��n$�f��m3nȠW��n�n4�`"Q�y�ٱIDTg �]�Rn�w�N{^�®��t6*��Vܴ�¾'��5( i�]^�+S���bq(l=&	l}�5�4���"��'�Dt�q2+�ݵ��XkLvoL ���F�.[KqL3�S�/�ki�7!��),^ U<Z+`�,+�+��R���Uvy��xU\��KSE8rE7u���A�Gu��F{��`�Z*.��H����e�iʗ��U�f ���=Lgla�b�e~L��S�p�_�����C/:���ۍ�vd��n *l�l��xcMň�/*����:�mhF��oC%��Q_�ƺJ�VF���A�!F�{lX��c�	Ȗi�)��������%m��u*���ñn�2h�5�K��U�E������D�ܯD<q�������Q��������ں�|���N����RO���[��s����3JŘ�4>e�A���ޕāC�����M=ۭ�7\���æ}�K*W<�����u�jt��A*���ژ�dY�8�鱗�HjyS�3>�{�ж}M[��΄��P�o�����Tp������wĞ���dӂ���wJ�$H[p�o�L��G�C�fKLal�]��l6+������e?��:Z3�W8���=�(���|lh�+
���}[�T����
�[���DFq'����6'����0[�j=��C�ZD�A����ꣴ�X���ӐZ����د�ȍ�k��P�
r�L<�.��	�vD7�I���b������l;F/�����7�љ���M�g��r�)��pHؚ��(�q�P"%o�?%S.��~'����9�ts�vPT�e�����I����X�Tsw�i�j�걚���+D6�o��%��U�%ex���ihS&�S����gآ��$I�K�b�~υ�# F�V	{.^*�
kz�߰צB�Al+�������4$�@Y�I��J�7ħo$�Ƈ޻mz�%��Py��4�y#S\���jk���U���'^n��n�J��� t7�غy��*x�^����uG�1�?��/���o�g�u���B�8��8nr�v�G�%ƆU��p1Z!4|c��W�!��Od�����
���H�t�� Dr<,�����_��uǕv}Oy[�5�}Fa '����ٴ������G�+�����*���<�aʓǽ��U?�y�����aE c�R�P����?��9x����Ȥy�5�r���7F���C6�:�jg�'�%0�M�� w���"~���9K���U��ZB�	�/�ƓL�8i�놞���X��ڸg���1(Z�B�x�nZ��?f�ʕ5�����ׄfNҒ�.xi�.4���:�C�*fg��[g�<׫"�re��w�j{��n��e�a�ߦw�<Ww�Q�?�G}}*�T�`K�s,W8��5QmS��H��"�C	�Z8E��]���2�}d��^R�/W�x������-�O,�c�jF��rgn�Y���`�&���%6�Y1�h·��±��KH��өB�ۗ=�:��w��-�NY(�(��\�����r��� ��!���/�5{�G$����sy���G�F�+�#aT���P�v�ON�ծ�x-����];�Wy��e�[�Q�6�<���i��Y2�QE��ݲ-��-�3�@r����ia0Tյ��넡��j���,p-]�a�5�B��df�-[H���I��Q ϑVg���*�|A�-ҩD%+Y/Jh���>:,@`�L� 0��Wpg�f=������L��{<�E5�KV& ]�=lĢ�.�β&#�|P������J�$��5�#�A���бShG���mP�E�|0ݠD���#�{�K;���`�o&�\�Ŏf��yݦ9u�=�I%� ��ȃā9���?C�q[�$����E��%uo���O�6^y�� � O
|�rr�N������� az��f'�u0�v|f㈯�5�(����S'ILq�fY�8d�H "5)����X��}ss@���1�k�[6���i�S~�`a��8��B9!�+�X�B�Pc�?o�G)e�L��U�3jd�+[g1��u�b�q��1�^=�	.��D.p��	��"�r@~���!S[��6X��-��rb�zm���+���`����
 �O��L�0��U��B({�POS�پ�j��I��X�v�2�UU��y�d$�X�����N
����n�_d:�j'�)A�ݡ,�O��^��ר�Pd?��� ���ݏ�mӖ,���n�$�YE� B�íE7�bӯ �a@k$��#��J�"H��tڞO+�<�k#�LPq��)/,���Qi ﵵ6�c/>@�W ��s7�k�z���m�qx��K�c5�E}����L��i{꩔#���Τ���>��-��ı�&�Wy�M4u���;�M�;��!7�5Xq��A�^�A^z2�.=�z��w2���,��E���X����E�˕V��l��~���c�8��H�d�?<��@Kͽ��t>6�N�x�o�ȭC�04��7r3�!f+`������}�(Z�1�F�t3d�4//j��w�6����6�A�����(����k{�y���pf4���~�
U9<�(�����!C�ZSVr֒��
ahD�1�m�α�^��O���/hBKY����6|��ưZ`D��hS���늠���Lg����^�=~�K��[BVx��w�n���o=wִ%�.�q��7k1��k]� i�}�&����h?eƷj�zV?�˙�zs��RG
��-Raf�@�7���qDk����#�Fۺ�w��M(e�붸���x�A��8��!�]v|����F�����0~חs��W ]%ڋ}K�6����o;Q��X��/��֐�CSo���Ip-jĘ���u�̥+^F�]QU�NI�1�Oq<�b��%r�~�%�T�i�{��&&Ԗ,���,��4VH��|�ѯ ��t���pD~�
�����Ӎgu@>��m�R�6gAn
�/A�'*�i�i���ʖN^����N��O�~��A(l�m�D�nY��m�Q�\��KJ��u�V�x������CE��Si8��S,��7'_����y��i��B~Fm�D����.eP)�_0�}u���3�E2���A����S�<sWC'����4�S��9��xa#��BK�.ww�����ߖ���"�/|�a{�Q۹R��.gS�.xn9�pDzmB>�<�\� �2��*�>v�4 �Hw�"�Y���|�oVlw�Ѵ_��i���o��koe{L>K�� P����v���Ӧ���w�dß%jđ�)�.(�$I}NA�2:>HC�I�%+zY���[�4�%,��5�ɣ����8<{g����qo&�ē��u����eiu=�����5�ڽ������xv��OP;$�,f��]3�[`K�h�n y-���;�&Dsc;��/�o�zׄ����i���-�=��*�+������x@>�?��Yq+c~�C�rO3�a;S��	}����?�� ����Ok�Te�0IX�v�WC" jM 4����J\��S�Rm` T�s��~�A�R��P������o�v��P�hhN17>JR]ւF ����޵��K�r�^���"=�+A���dv �1[�QW��o�i������YOK��w�%���+��t8��\����A�"��`���}��wr�(u=+�+z����&�ӭ�)���F��m�La}uhe !:�m�&pzA	��ߐ�������%�:D��m3-�]�#�;��۞;�E�'���)Se�[�v�q~�I3**����|o���@T��]>w%�	gE�`����	��0��-X�5
*���È[1��aUu��жY6C�">9@�Bs���>��(x7�Ҹ_�H��CHIY�}5�t�������~��DA͊���"�rOs�_�.\���o+�s�_�4V���ƽ�_���^ej��=R)����������\��/%�JS���2��PTM
���)˴�y�@��!�F�[5�$�G��j$�����7GOL��=߯L\��\w�8h8�|��p%��4�g�^�[�`!� N��i�1�i�M��qu����p%�Y�����ݶ�%h7Jx��L��� 9`����R���j����Ĭ����G����Fvܾ�"��4�Z�	��vd|CN�"��ng$�E7|�u�CS��n����wq����U�T�}��tW�1p�V�Ņ%N����[���0��&G�J`V��k';�5�����pu���]	�BTm�;Y�D($���[�Բ�Oͷߎ���/+*����
���x��]X"�~8^*�0��g�^1i���R��:fJ�G����:���5����]Z���Z/n�|LEO�ֺg�l�K��2]��������V�n7(-��U�c�b��h`Ln>Y��v=�f,�R�B�ĦQ��|U�ފ�����|A�S����WQv� �H�����kM���q�uAE�ons\�WM/��Q��7g4o��53�t?��=uN�C�M�����7�����JX�Uf�@s�h���ձ�_�r$���ἀ^H.=��~P��!���d���2�`U#�"(r��#Ӫ4��	�f�K}��(V�9/2!R�I��c�u#o��j�,i{GA�#d�\'ЎN?��:U�	�����2}�~8�����m��%�1�Ӟj ��h�u�󔺼hCۑ캶����7�-#����:�����2�u��ؑ��0)v�^�X��|k�N�7 RK=��p�?6Z_�(�����~����/�6*T_� C%=�A� ���TȀ�4��:��r��*��+H�1ˎ%���z����4���D��O������G(�T���i�^�%�^���M���ܥ^����{�dd
�KX�U旫yS�u�����~�y	��L����+H� [7��8w�]�p'�݄�78G���7���Q2{h<|d�z��ҕԐ�܁�Ui��\�eu�}��,I�d��Z����b�n���{��T�z ����o�~Q��W�-�Y�A�UT~b��b�z(�r�W��Ӆ�iO���(�W��H���Q�?�&�K0��z�T�	�qg��C�Q���!�ce�ζ���%⭸ᷙ�И]<����F�
��}��}a}�%;L4�\���|(Kb*�R��94-dH5K��3��9~+�$���wE�o?���{!��q-HXO��kX��s|x5�g�K�/N	�1���UJ$D	�Dg`���*�}Z�9�Jq-�r��r���=��i�r>	�PJ�t�S����]��k�h~b�:O�	��+�Rؾ����s�%��کU맸��8��X@����D��k���Yr7�֔�9k�p��ڗGyl���n�6E~������2EQ�EjM0g�"�����7Y�]��)��ci[��uE#.�5���tl:��U�K���L�N�-�db�x�<�rV�s��f�Dҥ9�3)'#����7�ה�%&���7�M�������n�;�M0�O��|�68�c����i����'�EH.5X�	�/�S�P8�6�=n� ��P��|�.ԗ����j�R�}�.Ŏ�����!d�aZ��ቈ�vb�e=�Ƃ�O!�0'��C�C��3� ����q���c~�C��Qfs\º:1��a����2�8���� ��s�6K'�����vK�����l���'P��G�����",
3�OJ>���#%��:�Ɠ�b6��Ŝ������T�ς�۾�y�� s�b���Aw�0�t�@��.��Ul�&1�r���6!�����Ψ�C�7�}4r�=��<�F} _M��S!P�j�|�F����Ύ��>����\��b�d���_�.���{��Zn
���X㵍�B$�H�]�h��j�i�Q��QS��ۺv2E]����xp�j�W��c�i���弃U9*]��f/��]J�<.H��'1�^�9Ę�mPܨ���T�z�Gnڄ �t���x�>��>nC�%ޖ��ړ���L��&Đ�ǎ����T���oN�{�$��3�U�9dI0X��0���r�
�T�$n��"Oޗ��{1D�V�
�Q���k����f�P�tBe���Vإ0.���������)��������V��Y�.��t��wHQ�Ӹt���!������p��W���� T�t�u�aJIA]7R�]�!V��n_�b�� A�Ts�8_�����K	���ղӝ���>M�u�e�3�������<�a�T�l{��F��Zb���n��v��4{%���]���@���I���z�~2m-=$o:��8Q�F�5?������"5g~;q�V�}4Ì>ά��ڸ�Բ�o�� �r)b}ɺ)�%�9E��WF�?X�/��"��mwr�M����� ��-�J�ʮtL�E,���d�1(0c���^�w�Q��O��KjŅ
RB\~ڋYq��)��� ��Tn.��Uy�VD1�į����y��%'�\3,f=��4ץ���Bʈ�>��^��x$~��3H1��[H`;v#��s��o����~Z����J���X�-d>����O�&�{D��	Z��&�Im�K�A^�P�k��GVdHdA�1��;����E��8B%*��>I�8<-�k�-����Ҟ@�F��k���{�X��5nG�p<�l��雷��㝳�T��r��{���%Df8�ƂY�F��""�^@��a1���T�o�+eA�D����l�M��Ƹ�]��3��Ej�z4z���&O���c�}���S�� ��3�R1��$�b��tn�LU�:��3�ZO�%��>T':׭�'q;�|_����:IgB:�Ӧ���q{�i� ��c�fk��KD��-�ZFZ���L���h;��нi����� 3�g�Otg�Uc��2���t_���3�p<�Y~��z���6oM	���1D�75�ٻ��.	�:�!�������~B�DG�.����;M�g/������0�\w]A*Pc'#+闒�
<�x7��8pC$�$��;�Z~�z�{G
plKi&#j���	���c�>$ݽ�ˠ�1v��?2���
0k��L ������#�y�g�G��I�%�B��d.x�0��z>�'�y�S��;P�J��E�R�\�����mÕ��^�#�a�������r��m������O���ߵ���W9���	5.hI���g���#� |���k�t�獏�2�;yw��Z�,L�|��iJb��%lуp�.���IgzC�0>,M.�v�t}�yDg�l!]���p�qHϯ�k����|>n�楼�{T�t��־S�6�m�PZ�;Fg�戔s�ĞGz���-�1�%KY�@f�qr �F����rR��$(���8���O����,aF��  �X����6�~�C�AJT����8�C� �7{O��pj]\=��6��$GV �=����u�VT�:��#�KJչ��'��`��
ّ'���
�2�2�5���G�%Y�B��]��,�s�/Y|�8k��Z:�<%g���nP�����
�ß���	y[�<���t��0���6���ˍ�T��:ɓ��&�j ]��UiLHG���p�y&�D{�����$�N➋.g�f�a�
u���w�B��F�s��e@�AC�q��wb�	����wR�58�}4�ءˀ�e��������qȻ3A�g+���o�Ph��n_+�_��߽�$Je��Ag��BO�m���$�[8�1.jC��3������W��� ���@�ʽ�G���m-��F3B�a���ݩBkM^��YA;�����͞UIjW�k������U�$�z���6��]&PG5iE��3pz�&��$`� g�P!��k=%���;�:���!2�������6+�fP.=Ѯ�
�0Dч|���9�v����Y�X[��9/ٶ��Z -m[1W��]���j��{�u�)m�� ?��7�j4t\��K���x�M�+2��E�T�gd�Mh [7�%���>�zS����QsFx���5��ȧ3V���z��;�(TI+���枡��PR�
�%��]��{�����6�']�'��^�K��K��hf�Qၓ��aW�/��*#�i���	�e��،M_j4�)�u^j"�iM���E
��ڇ)�[R-Oc��S�� T������u��p`A#F�-�glW�r���4�d��ؾ��r)_������,/.�S�]�	p{$g)쮭FUw
]|1�VʧW��5:�ۙ�s<�̔�Z�eړ����o|v
a��fH8�7��xU<q�Q|fa�lX�b�N���9|��_D�V�w��q`�$�ڼD�5�e�1���+���rj��3����P���W:ш�.�b(d�d}��rKZ�0�S������|��Adگ��Η�&�e�EnOX��O~r��9�	s��(�4�;	h��/3%�e����,�O��8d������� �_�:�u*��]���AXhp�`�^ַ�%�4{w���|�=�b��Wm/_�_A��Ҁ�� ��(�g꿩Mi3~ �K�>�.�Krϻq�k�����'���RpW�p�W�����j�hp���8�(�'�e��y]����kf�����e�4<�������5���wq�o!�3'`b#AG�9E$��GgN`���Z�M��4�~�&]h�-p�7���fݘ�ҩ��tk��^�Э�҈<ٞaBFK+��|4LÊ��K�+;w%BS�d��F���T_�@�2LR~��r���f�_0��]'} ��i�m�:�"Tt"o�XI���9;��������{�}&漡1��D���HY��1�ëI���EJy� [&���aN����w��y�����҇��J�L�ӯd��<z�3�����>t�L�akǭ�:  �����m�Ti��*djC���x̐���D�j�'�פ�����wu���'$�<�9���E��c0���6��.<�f���'��4x�v��F�u�	���х2	��^�yC�pԙ������-8�����Q��L�vj�GY�`N>�y^i�:ݜ�h<�&G�ޯ�b���\�Z>6bI��e��?6dg(%�x&z}�x�Γy�3�Z�TG���4	TA���׊�oT� G�o�+�Z!����M�������4��bgAJ�)Vd�  ����]j�2�|C$*��=�>f�U��K4���`|XlxVHYEB    fa00     8e0x��1\�)e�����tS��I��C~
0���u�t?����~b}�k�c���m�;���$8�+Ex��71��`1�]�Ñt=���&�_Э����3E�E��8�4��U�Ᏻt��z��ˈ�
I�ِ6�l���E_�!���.m�P��:�3�a��5J�5!%>��aE�{���9�����ClR����`�J�pzb�w78�~�j���H�I�;S�bH�4�Ҭ�V��=��	������S���pO�� ��(Oͧa,}���v4j�������ſ�a�!ri�m��h��jxj���)MP�t���F6� ov�h�ǁl�d,��wKp˴�]S��*fǤ£N�"j��N`�e���M�Zz�3Z�3��V�d/
s����4�-�.6��A�e#4�`x��@�������i/�Q��#�E�i�����U����ָ�~g���w��0̮+q&B�����Y��GM#�2j�u:LU�C�1{�P�kˎ���mAM��u�ҕ2������>~�&���A;�v_��/\0�+�<Ah�xQ��)���!��s3�&�y��$�[	g�n���eNy��]^����нopa女���z[��4����y�"!J��p�.�0����LN�z�o[&�/R�o���-�A�"�aZ�:�I���Y���tt{���BGwc��U ���p��Q*'�6}�j�ȳ/�rW������}o2^�����J����2QT�i�e�m!.�\ܨ]TGj��d#]K�L"X_(35\a8�K9���[�	��9tsZ��и��HAz����M�u�E�bn�e���e�3=�tۮTud������lN���
НȜ�������RW�D7LdA��l���/��}dotc���\��VV�s«;�Q����r U�v��@����U����Dg�F�$Ӯ��t�.��qd2�PM��;7��cA���g�{I���5R��X�(%Dv���8Y>�UW��l>C>	q*�,�8���b���}k�Q2 d0�`�K��)�������"/RgGt=|�(HP�#��P1HLp�����4L�-������)j#!c���?�
k�1OA�ۻ�
:�1�Ov<��5�< *�T�S�ƥ;��f��R�,i�1�4��6���ܜ�����oXR	��	k.����U�3��M�L�����榼!����Щ/�w»�~�=�7C{��f�����'�$	y����C~	_��.`?h!0���=���+J͞yjo2����3��8Z��C��z9�_���|y9֑4@Db.�:5?�Ү)�c'��`*[�I_���݊l����@���U0��:3�_�m�qH��G*���8��y�Z`� �Q,� �2
s�R'��x,�px r!���ٯ<hRRP�_��^th��X�_�Ң�cɯS��E
Sč�l��]�����G[Jc�r�ՃL�>�xP\�W9�U��B��J�`Fwam������j[P�������U@�����D�D�����'L���	i�� ~�0���2R@ b���s1��f*�QΗ��IZ��yx"v`,� �ɡठ�?y�Zl,x&��ë�R�t���n��k@V�k�px�ǯ�پ���ΈOɹ�����+x;tg.��@��as@�f@
��mv�7E�d�Эj�^g눃#G5]A��@�:�XB�^�~d W.�pn�3��l^���jˑ�j웎�IZ�M�	Ep�+�����_z3��9�}*��i�8�u�	A>$����4j�uvs�h[:�kN��~�_�ȯƊ�*`�z}"��βĚ�H:Y�R<ϱ�[}F�6�W���$�~5�6���k�n1F�� !��\W=#���<C�=��-lP\���&�}�R�9;h�V�T1ٰ���\> �kT�qiU�?)���Q�р��n>�mcX��]���[�$�q6��6+@E$cz�O3P�5�Ś-���I��~��Z���	��c��Kr�l����;�f�Rd��3�p����6�,,���]�	�'���1/��R8V�9�v������zi"�8�*]�":C\.��8�	!��0��vh� �-�g��%;޽M���L�_w �On��YQ�ӡ}�$tZ���X��$f�IK	�aXE��4A���[��YNZX/8*2N{sE��n_��1a���$����%X�(�6�n�a;�ԅe$�i �� �8([R�XlxVHYEB    fa00    1110G�|�����g��!uyf��'�ܚװoP8vtr�{�*X��-�y���.�#�5g�����Ԡ޶C��	ˁ/�ɄZ.����^+\�d�bR���-�#�@4\�w�x�Y1\}P1'�z�>g��b��iiω���I�� ��Zu_�|`(?S��~�Q��V#�4* ���Vp&.��_CID�^4�{�o���"u*ܘj�����x&��7`�q�Pn��XÁ�D��X.��+"&��o*�z�D��=`0:z�gΜ��3'P�����gf���"@�	x%m��.����㧬�g���$Y��d�����w��9����-�9��[1�Hd
�]�՚�(�%יxd�v�ъ�C���7�R��9`P��	��|ҞO�b&&1/.�2K�N���+��/�N������n�3 �ȃ��R�@��c&�:>>�g��u
:����WL��[T�|v��	
'b	1�g˧��H$��8�/Z�V82���!��
�}Z���Piv�޴Ҡ>�6�k��SN5��*���!�O�C�О�t�).�"����%�V␋���O�@<���˅hkC�	S��3�%�!�ܣ��{1Vd�kSơM�K9'T�Z>x	YQ��l #3h��ԏe�s����]���R�_di��S��X>,�s��Nj0����I|����٢#���kx�����ԕ�M{�O���X��j���������C�b�4@�p$%��i�*�����Eod��1��l���M�`T���4�ӆ�O�R�B�[rx��G�y�O����+&@u���u~��� ��"�`����s�K�@!�(��d#lR����99B;�Z+�M�����fw�]�����6uTc��v*��g��tۤ���RtF��4�Z���8g�U������O�"0�7'�����_O��J'����(�!�y���V�13��H�-L��6����i�<�� M�,���Gu��� �:�/�t��[�E��%y^`a!�e��F�T����s�*����r��DN����w׊?H�S�2�.����K�B8��il�\���Ҽ5�T�#:�_hډ�r���Dn���KT:E���w-��Z�Wli %;��i���(;�O#�+ ��{:��H`��m�3d�;8��������x̑P����Ϣ,�_~��X�%eI�ԫ�G{`�AC�1�&�s8�gɡ�wa����Z����C��B���7�S������cE�Zu��r-���}��/�C �}�^�1 ���J^o殆lLȕ!V�'m^h8l��2{��혟�n���
��l�>;e��Ɇ��f
f����êE�Xvk��_p%�@rB��E�G�<+2�f��{u��	B�G=����6h�D�\1uZ ��JZ$���td�5f��g����^*>�x���hygQ��&s���*�X6=��������N~&W 8I�: aQ6N��G���7�i�,TyS -R�EO�e7���)`�N�izXҕ#�O�)��?�C�"�ċ��Z{Z��R9�����:��
�WV�>x�9�H}�����10a�����y9��N�[^�nn��Wj��M��+�.���S'�}���M2��7�U�`׶��)_(���@p���a}=�������;�>��@�F��E�$�yFe�G�G5G7[M�A .�3{:�ʯy��A_�gn�X�q���$|иl:X֘��I����7z�^�i�5��u��䑛?TI����)�+5�t��Z�6�ל�2)�^,����/��!�SmM.��V_(t�}��_>�ue���>v�c�7�O�
7+�_f��ｶĂ�)V��Ybl��}R�������H���`e�s|���W�ʃi����eu;��
�Zac|������um�����t*�n�`7'��X%��~d����)�m�L� .u�D�?R����$��N��ŗͳ��Zh�L��b���Β��^��M\��'rYa�ȃ��Ɣ��.��GUZ���q�����@�͆�O��Zn㞅 Q\�y����<�_.���H�H��u6xcÐ�S��=ph*�܀r5���u�Ƽq��[M�9��%
CQU%���%���qQ�)J�7��G����{���v~��왽^I����خ~�&��#�#�ib�ٔ��+[6t���r.H��Zg������K�Wtݐ��j�d ��k A�$HA�x��}�>�%�Z����wE��A�B�����z�^�������8��}��G�:vb����9,t�1���1��m}��]g�C��]����D�[?���.�;�
c����*������6��R� ���/��?�Ie�O��ܵ:S
si�<���n%2
;gm���`*�B�J(�?�@��I{m�:N�!����I���0x�"�3�q���S�q@�Y�������(>=������O�&-Is3���B�]9�ya�)��A�t{�c�\1>�w��P�WQ�a0�������Ʉ],;Vvf,k.�)��3�!�u9�Nm���ԃ��>0�P���r��Xet	�fG��gh�5V*�ǎb�AJϲ��#\�|��Љ�֗b|�91��.�\,�n_S�2D���h,p))�&��C��y�o���� �P˯I.I��&�=�9������HD?���Wi����U�,��J58T�
�h���i���TJl@פw]qbN�n�=�p8���F)K�'�N���s$���.a�M��Fi$����"�)���B]a���$%�F]��[���:tz]����̻꽢s$��:"GܚDhרnrQ�:`�;0�!�.�`�ӱPȒ��4M[2���X2���g�wh�=X������z�j��fœ�	h����v�.�ltY>n��غGbߦ>�2�}�����b���B�C��0�M�A/�o��e>�0˼1��[� >���D�v�1�'�1O)S���>N� �-P���p��5����5���y���B!�m��$?8��I'�?���3Q~N:�Pl��޺6����k�n�Cv����	�;6��tZ��d�V�C��e9�� �O�>�U������+����)M8l�휉{@�jZ��ǯn���߸��Ɔ�QZ�Sڣ��?���T��7��
�ȅUIv��q:�eШ�$�$�7�d��m�7��wfZX�ϲ�k����a��u�ζ��;���(�4��}
2���շy�������h��P�
D�}�lhR�y_O�<U򑆱p8Ǖpc�ܴ�7��Ĥ���~<�?�?�-<M���F��K���P�:�{�	� {l�3U,K�n���T`��pK!��q&w���»�`��~��x����M~��4V<'�w��9Ǳ����˨���L�=S�Xg�h҂����"4Y�je�:�8^W^mkF��^�����k��� `{A�ց:vDvW^�gV����u��0�9���6��Ѐ��. p��
�wj�j�(M��OI���SKt�9@󂭅P��^%�5Bـ�v�ᯗ�ř<�=�97��z1+�o�F8�D}SI�2�`��R��~N��F��ʁ��.�3^{}�()~�����y-{N�7y�k��'.^�I�o�`+
���lk��e��s*ڐ+0x0���Y��:�,�V��J6x����3B��ƌYZ\���>�g�ɒ��L������{�أ��_��=�#��yX�k\j�����dhs-�ȅ�*�2�C�ր�vf�?EV��xM��5OXgΏF�msp�~�w�onb��rRN��e� ��Oyi��Q��~�6er��@�YH�T���T",��Z2XWD����1�����,\6G4��\�k۹G�p��ǚ��hE����)�y������z��uM6�;}�)����MZ�V���� S4�3��Nlc�Z�Qn��ر��w�V�$0�n��߄v�#�^vtW#k�m�o5��m�|]]pV����^���.}wc����c��;z/pi]�f��p��"��?lf�ߗs4�oD�u4����ƅ=�#>̏|'��ug8�p"~8*x۲#X.'�@�D^Y��"�2v�r�K�j�Z�8�#�ūe% ��/�� ��)�����8N�ҌXR�+�.��MM��=�X���0©��v�=q���e �����c�˨��V�.���ښZ�O{�����?Dn�hG#FɄ�<QE�h	������؛C�.GuEH�>���þ�D�bxG��ը��vy�aDᵽ�6�XlxVHYEB    fa00     ca0�W<�"�����x/�S�ȩ	G ��-d��	��'P�(�m�2@��h�͍�d����{)�������6%���/�w�=g�Jf,]\�Fn�W�m�Tw�11GO�L�I[�U �V��K�(G"�0�qs'u�y��������|f�g]�W�ڸ���U�oXO�P:�ԼH<�o7����1���%q�k���$]n��\�*����~�1���!]��hωx!����0�����$��00�C)ʬ�!+�U���������R�_%��6�� -Sj-EZ�f����"!`G�g 7
LXp����[�WJ����,2Xg'8d�-��H�٩f�fX*��O���j��j�}f!h�s��"s��*L7\%Q_��Z$^�e�p�K�֡�1�%K�K����F�eOMx¢K�-�B;3�iժI	GT�C��|a-) �I�O�-.Lm$`�M> f��%� �{�S�9E�DR����t=OVgh�0M� �)�G��n�M�u�����n�^qg�x�<����"�P���9����:�kKN�VK7y��z����U�F���H.,3���%��A@�v�(L2�sƔh,�^�aw�C�����rב���>����A���O1`�����tbQLX+ĺN��G�P��oڗ���Me;�gV�(�m�V�t�uM��U�=��Q�(����`x���69Y��P:#��7MDe$�(�#��M%�ł�>���<�̂��~���I�y��IHg���f!ԨC�(�	@��
J\���00n�Y����z�.�zR���Q�K[�!� 5d4s���:�9��{�W�X����\h�&�	:#�3��i��kv���B@���6��-��TqlIf���]s
��z�?DB���a�J���n��}��L[@Q�q�Ͱ�m��%���X�>��*�FD��)�	�J�����/K@(�	��&����ƽ�= ��Z��A����TS�����^#p�2��y�F�+�3�J�2�Ì.xw��=�m���R-RŦ�s`6�g�#ť��6ĿI13��K�s�v����8���{�Q��ꍮ�.Q�ƚ�g�܇#��F��=X���J��WS����*M�0�my_V޷���R�!%�υi��&oB	z(�[��O= %�7y����^���Ë	��_n��d_}H�ܶ�T��z_�2��
���i\�[% �����г��;�y�������'
/�^�R�d̻��/�7R�}@���\�jTҞԧ�`�\�d��`�2^��g���������`1�������}t@al�/`c#�:�	�����EV���'1 >,�	Q���j퍦_qi�^c����Z�޲����z:�
�߯� Tj���8?C�q��|0��gV��(W��2::?��<v06���~Ӕؖ�L����|j/���G�*)I�v[X���Ɨb��^�@����͕�"x���e<R�~��q6P�w�L��D�pO�^sYYf'>�~0�92����p�s0�����}�2��х�2|�,��A'���\���U�K�b��"��4���I�����$!*�"tA���W�>�x��(�WOZ��R�_v5R5�_�8��)�n�t�?֒7%�Dʔ}'K������'���%Hi�Q^.E
��Q��JF6��Ƀ��+�/�V}�3lX��%�[�b���h�����VZ|4Q�H�(Q]%�}���tD{=��
�e�^.�I�"��$<�O�X�X-�L]k�\0"�:!�p�	ֹH(�6��,Whן�m�������5cR��t�Z�oIǖl�JP��mr�(�UuC���&�¦?�2����U��+�Tk���דbߋ�5�v�X4՘��&�BԵ��t�,<{���G�\8ҹ�����YCUx�0l�؎=�+�y�QU^�8��N�6H���v��^��$�8{��ﰣ��
վ�'*�{� /wx�zj1y�ng���v�KɄ�
3Ҭ2��m�ahT����Up{e�~��~��׵m?�`�|@�P��eH��$2&��#�ߚ�6s�-�? ���?�O�Eh%��D��;$����Lߞ�~:!A�V���6�F�ÐD��a�o���O3����o/�e!�q0 #���X���dK�h/~�O�4#),����B*^k,�E�W����R�"U��C¸
Ô��^P�?:����@ψ孳�	���YEv����C���{��Ө�"�,"CW�+�U�A8v�3�1�A*O�r;>ƈ�_">�Y�u;reNtRFL���KF�A�
�`ƪ���i<��C�����	��|]�?рW�6�WP�wƼ�p;@.�C����*����2�����L\ۢ �ŢK�ǼŐ�ì/���iJ�ͳ��������|V��BmW��.k�o�^@�~m��?���Y,��j�nF����LA�s|�w�p1U�ޚ��my���AG�a�)�Emh��0��Sމ䥌�\�寊�6�Ǿu4�97�9�r�L�p:�95[k��<u��#"Ӆ����؇�I���N����}�s$�2`E���R��)`��`�����T��:oӜ�vlmb�l6!�8cMz�+SRt��P-�� N��v
)ӊCQ��xf�%�x�$tj�1�+��Pp�,�E�ꀭ�y: V}>��%8*:���e*Z��X�Ѽ�JK���� �z�sYe�����[��yu��U���R1z��U���?P  9���%��wb�q}5m��"����E�kT��y��L�J��LVO]����)<����땕��=o=�����}q��;�����IV��C���y�ND���,	���8J�Z��2�_+������8�%bӨ֘kn�DA�/.wP��$���4EA���)�p�u��1z�IU����jv�0�H���������B��+�]1+��=?khN ��f��{�����Ar@��-�RC�y��Ic�[�[�u)]|���AD�na�W�C[���lyf��t ����p�o�Z|��0���C���� ��Y���k?��6i���vaz�y:�k?%}dp|�:�p޵�T"wFwT����{���_٨�T���g#z��y�������*G�O�}���n#�H7�Z�/Ҭ����L\�>��n��{���V�XlxVHYEB    fa00     3f0�5;u��������n��7�#���X�/	��?l����� I_�n�g�b�(?��,`���o�)�����n�x�7�ۆ�9�l!ʖX���T��V±2��OJYcčI���!�.�ԼY~���2ͬ�{@L��y���G���PGQ}g�U/S��}|�9�HI�nX�JaPy�i�	���ƅ�&:(EGvYU�^2�eo�nMCBě�S���E�]��:�Vw�Hb9��NmATF^d����:���sV@�$�{�s]�
w�_K�����x΂��q>H��CKY�Î�n��o��XF������Mn���Hͤ4n�V�YPiȑTV{�(�MO,�U�h�Ʒ1�Cy#������/G
����)�������Y8v�����(�8[�/� u�%(��녮��~7d2��K2 �Y�Ŋ5BH"ߠq��dH�qv�Nm�u�>��T�ҋ:�,��:ʌ���������aE�'��G���Bϥs��_]?�uCYr�pLEqA���N�C�Һ_@�"#��ƲQ��҉�g��j"c&���'�e��gel�ʿ����)��[�D�ĞT��m�y=������������N��`K@�=�zyV80w�y)}iA�Ai�_:�ޣ�;��j9��՜Ll��[�l:,KYs�z�B}�M��p��6���Ӛ��t8��W�����̾��ۜ��o���0a�9��ye-U�J�Dܷڦf4t��.d�'��w��7��R���)��.���5������j֍�pK�յ(�\s��)n Z�Vg�����[�� ��AU�����:D$EOq�	O��+O��ӲǷ :����N#vwܤ|�ҫ���&\gZ"|䰎e9���I;ߴ��׻�>�Q��y�u��	-�,�Y��]�M[R6.g>�c�H���Q�*o@]��9�7v�%x��q�(�0��:�qR��PBl�`��&�����~,|k�\9[�������	$�}����{j���XlxVHYEB    8096     b20�Ʀ� #h+
��pm���}? ���<�{bFOB����Ѕ�q~���'��-7k�W�$�u��%z�C����`y3z���QkC��XO�U��)�6\8���'��۞��93�]���n.�D@��xaZ22��0���TV' ���5�;`���Ǹ�����7EC�n��R�@��v4o�#��ғ����Z�j��0">�����G��@���C��m��9S9�*YL�e�.�����`��Ph쯿d!|��h�:����v��r��t�"�9�#�G�Ze���z��I�H}��Bȴ�ɢ�[�l|��D����Å��ԋ2z�_�mR����w��3��a΍���(G���r
���O+�qmd2�*�a�x12Ulc,X�]�g�Kh��)L��dU�dE?�f�%�%�L �+��(�d5��K�4��L��G�f�i�t��R�� l�D�I*�4�v�_Lױ�e8�p�~�Z�CL_N�s�=c��|�P�@�	��J<9[a)@H�0fX��~�v[�����2��>:�Ƀ=m:31��}T�J�w�G�i�,�Q?͛�N�Q�Xq�� ƨ
��Z	���ƥ�Գ�6L�"����>�7�W��!Q.��i�T�����Xoz/a2i�r�E�X��R�2֨��5뷧�mq}F w!�2p��v�O�/(�,�^�����3�c�`Kw�4�0nrx�b�����kq��۲��Q*7���n5��2e�K,��*V$���;��ٌ�,����i�,�}�D�����.�EˁB�(��%�X��J7����=�ˑ~.�@����sH18�(�A�����ސ���5@���۰6��w��n�V����h}h�|�����J0CY"�;������0�L���~�� >�~t$�3k%4�1/T>y����;�s��2�I�=B����X���c�DGo.L��	x�"��x�A��Ԗ�4?�?x���'  V�D?�ʴ�ũ�*G��a�6�Qp=o��LJ���xwOODẞD�D�+�auf�֮ӕ�i�����Q���˓,�A��q���%#���T`�$�(�E��p냣�������Ӫ5gshy%
*��=Xhd޼������W�+��5� u\&�}�;������h�J<��*��'!C����3�Ji��D:o}$B��Mo�Za@�s&�F�1�&
{����S���5�)�+���T�%Yl�P'�h�t��]��׼x��Zo���X�c=�'J�L�xn7-n�3���BG2?��b-��J��~����}�w7t���DFt6!H����x�o�XƐ��t	�թ��~�#6����wϲ���6�S�W�pp��#x�:)gad .x�#��ϫH�Í���TO������]c�%$ݹ]T�I1/�I�����HXn�VO�������A������=]͂*��:�T>�D����}����s�{�ø[�y�П��q��s�S�$�Ԣ�+""	_���L��_��N+@'0��b.�ϫ�)�S�M/��{�NP�B^%R���<j5�$�z�0`z�)����c,����:���Z�@��d��q����M�0kJb�ʽrV��ܐ�*u_��C�\VG�'h}����T�u`��S�r�A$���>r��-e�cF*�\��2���ج�Ջou�=)�&t�J�͈�~x)��J������-��]q0
�5k��$�q	�U������	��g:؏f�_���_���)��~bG�,�0��M	�(g]z�ƙk_���KS���{��3��CG���&=���A��"Cl�wK�T�ƣk���Wߺ�^5o�:#
��/PR�@C�)���\)v�{>�7%A��*?A3{�z�5���1�٤S�W�1���>��uX&�Du��*��޿f#_fAe�K�1Fd8j4�	 �KP��sΥǫ�/l�'�����ڍ��8 >�+njɒ�ٴ�-x�\��_�i']w*��c����z3�C|RB���y��u,+��쇁���#JW������c�mD��AIr
�Yf��`e)�%1�/�f�(���Fn����L�|�A���cE��$�&n��.�M�8L�sJa0$�نĨ\j�����1!-&���S}��_��Dn�����j�����:g�.XmW�ծ�$i��e-s@
�u塷�X�O,�'�=�}@��[,-��.���S�o8�Φ���׽�k~��B�������������m��t��a�X��ZZ<��zp@�pl�"�I�ePÌ�b� �a*�ױ�ͼ� ��|�t%
���S�vl!l�O�����ĮZ�9g[�� �/�������g�Fᆃcb�)�xYD��)I%i��KQ�v����u���Ͷ��Š������>����0:��6��|] ��~3�Nus�������hH(1¤����d�Ԋ��<$Ү���]���צ7b�J8��X��"Md���E�G�UT����n�#�O��<�K>o�
H^c����D#�R�G�DZA>'���	��
����4� �
�b�ǭE\�׸�er����D�0�p�m3mz!|����������w~���y�-���L�)�"��%}��pC�
	�\��P��L�Lx���"/�W���e.Q\�H��uю���8M������s{��m/n�.J���6�Lm�"��˿�-%a�>��Y�#��k���-��ސ�,� �F��t����F���t�*edV�
L���v��2Ĉ���=���`�*F���Ó�	��q���ੂ�@}g���oI�ĭ�>\}I����W�%/4�