XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��	7��:4�e����G ��r�%�.I����a`7��#���l�y���hl_C(�"[+�W���ԫ����2r���Pxƺ���ӽ�ݼ��+�«9�D
��9g;d�Q����0VUʢ��F�~���7
��TRz컓3�c����I��(���A��L�#�������Բ`f[�-R�"�A�®N5Ymt���=,o㸚/�S�Qrؚ�6����#��v��u�rp�Fiڸ@ǧ�j�Sd�q���⋁�u�ùek�J�i�����c;�>�O_�LI��\��I���j�(���V�b�=����.Ah��<�;�2��1^k�|4�ꎃ���itp�bʴm���I%o(�]�H�[{�5�X����v� ���"_��
�c3���j-�j�U���jW����K&#�tH1����,o?p�ѳ?�ȣ����lJ��8�0p�KV�w�a���m	[ݪ���8�B@�n�a���ɥ�� յ�f#+B�'��7G�
�;߻��z���l1E�
R5`�6�3��^L�U)�L�'�ͣ�Һ�0�����W�?��V.u[�{��@&9�F֪gyPà-,���bc�i0�m *{��Ji gP!�G�Z]��������"h?�����q�x��6�hw��^%�uy^��L�
I���
����j8%�X�2>�����)�ۦ����G&���7N�������=�O��s�=�>��N�H�h�^�#��ͯJ����QC���4�K&(&	��㾄[x%�d�&%T��z�XlxVHYEB    fa00    2040�/zk�<�9&V��o�P�;T�&&̝;J�ie�M�t�`�"�����w��;Ka�7�zlcK�eX�uP��ű��d$�9H��g��E�y�ք ��/��g̝��_mu5v��L�[�����>P�ow�D�`��MS�ŋ>��5Lq7�J8e�UWv����:��}�q�`�Z�ߦ���ѥ�����Y(wq��������z�8%��0�����}��a��Ӷ�����"�M�=r�Nb<E U,�S�_h�љcd3嘹�|�*%��Zp]:�����=e���/��;���r�R� ��3>�T�9��9Y<PV���54�0Ue#����C�G-i��9����A���h�D W6��j:U�!�;j�lݸQ���'i�S�c�~4�#	$*p��Y�ъ�Z��1Tu6�;6ںjo��qW�X` 2Y6u Q���]9�2d�ue��@UB��<qR�+��r�V"{��WKByh��gR<
�-p��kt+h#'f>!��H���*�ݨO�|<���y���I����yiq���ɱ����e�}O[�Z�$���*�TBm[��q�f�VO8�bz)��K�<u�&y��0��QZ�/�Wj�{@y'����\���h����k�v��S3��rԗ����r���H�ŏ���}z��߮��)��1���c�{l��$_YoV[Բ'����#QC�n�(X.��P��]V;p��|�t��G�WEނRۊ��Hw��X��鴒nR>J`'>>�!)�����Ưm@,�*-0(���7���mk[蕐���,G�G�L{b?�*�W7��3f*��� ��sbנ���kC��'�jv@A�\' �iI}����w��w��}�AQ
9z��(Fh@��71�����|l2B�1l��8õ�I��pWi��p4rt��u��[����1�#p1����^�Ke��b9G�	G������ߤ#��	X�ؤ���j�%�����ilN,q�w\��Y��Fz=�dW"�	����pkX|��@)خ|VSw����,ր:�h��(�d\��	�Е�z�i~�IL%�O��G�Fr��7iu����D�0�Cc�1~���xЧ�|�*B,uǆ���ָ$L��3s�*!f����eBqRHm�O���}Lex�����s�/x��颮X��Ml�������y���O��
1����u)q[fN�Gi��'�l�?�d�t����?.#�k����'�T��ۖ�&�)ߤ}�mw�q�n9�xT����}�x�nq@v�4s�3C*jt�{*�駋w�h�ܓ] ���M�-�3z�U��}��md�����k���ur�CL.������6�e ��Z�l����e{�ːY��d�y iU5Q|��� ?ȇ�PgOAH %� ���l�d�D�J��8v�<����(��xӕ?��EBl�4���V���`8�k��Ҥ�n�zpKjI���R��<e4��@#��H井y�1�Tf��m=��7K1��M�f�V=zi:5����tɎ�٘��s��U������zFÏH]a<�뮞������X"�S���d����\�;�:���n�Yuy��\�d������� ��r���a��{�Ղđ�F�v\���mR�gд6ɨv��|K�������j�����'��&O��%$VO�}P�wayS��D�m�-'�][��B��������@n ���l �Ю��cJ����Fҍ@'8=-�8�q�=*��x��'g̫$��f<d�K�6%�=�$�C굿�T_�*Y�(<3��^��wr�O�G?�ꎣ$~!�5�n�d�b�=e9Y����S�\Z�{�^��R���SIk�P����9�ph �N�i�m�#�6s�}�0U�9���$��C�'�^������c�!�%��v�1�IYγ_�*Ry���w��B���#+~
;�ˌC��%Bb��_��ED���-�V�s��I�_����&o�u�?SY�3���R��2�`��a� �Q�%�8|�a��Y�R	�އ@+5�@�"���&����koq[����W3@�?��ң��Һ2G��ӦԂ%DX�~��4���V4�n��s�l�?�����85���ӏ��,�=�;`�{>k뉒�w� �P�F�~�V�ZK3���g?̟��x" �R�[��|��x�_yM�Y�88���5��|M��۫��#L7c�'�v��L(��!̬<�Y����e.��D��IE�K/2�����	�)EW��z�J~���t.i�ޅNA�Q�係ϔ��?=z鹊ɠR偌��R���3���b��X�E(�q���2Y~�9"P�3���_O��H�b�0S�����8*��%N�8|D�5:B(C^�@>A�v^$��KBIf%1�%ਟ��P�?A��b��w�n�F����6zȼ}1h��.C�G�3P;�q�����K�. �^Z����b���70d9!�NA� ��;���b�I8��~_�|�`�;ğ���9�Of\_m�pz^=q=�����'�W����$�����;u�r�:��Z�\�uW��ѻ������͆��j��R�枑Y�o:�!��)��%$c�]�6��/_x�`y�=�LE�����c�9Ŕ1�	�fu�(ev�/�<���y��IW ���*�͆��_7��ᒄ��z�V�F��P�4��M��[U\f�e���&|�IH�Q҉ːB==�y9^��#/>߅������!�Z{��D֮�����(r�,ӛ,�Bs����`bq&0�b�R��1��7�%���
J�#$m��O�*\���Qq?Y��x�֡�p���[��3 �`r	7N���W¹H*:H��XR3�_��2���CU�:?��!/�Յțu�f�8�Y�E�1t�l�+�:���蹴:��+��c���*�qmKt�����;Z�x><�C��&�|��d��tsd����5�8�A$�M�7�y���%R�HU�	`�
4 Y M��p���\���J	xꥢ�iXT�L������T!���>A���^	ϷY煆e�J�"X;�Ƈ�8S��P���)��g�C���.PV�_�G�e����s<��m��^מ
�1�N����&.�ǩd'���p��+7�9t�UDɖ5�H�;��i3.�Ϲ����bh4ܭ����,�&��X�>;Q���w�^iAlʗWm�S)�U~���bK�K_S�ވ���C���E\�Z}�Mvs=;�89�~����p��_����Z�7 ��Z�����<*�Pٯ�,��Ӥu���@�ˮ�d��[�Zݴ���iq�4��B���:��`��`�0'ї����/؃>��j���8"0�g��im�qf��$Kx���A��3x��_"nP!�y��c�8�etȱ�9[��ٹeŴ�9Ѧ�ͬ��^�>1o�p4ʍ�FX�@U #��f��&%��T�	h�s�ݵ'Vۡ�T�����H��UE��E�PE�����&>���L�ІR[���
��r�����uKH���u��܌M�p��E!s��τ
TPv$�M���e�)�>J��mN�?�Z$�Ŗ���y�v�Ɣ���}��x�B$�Q'���0Gg�+�dR�*��]v�;,���� n���5�V�~z��D@�6�궞o��&�ޯ2
���w�25������t�	�38����ۧ�cm��;d�1�@ץيw����g� |�@��"�=[���"�<��d\�1b�Y��uY���R����V>J*��
��/W#<9Y����߹���U���d��p�"���Y���u�\m/R�Au$�3�ю��]q�w4 ��ZS��a�U=cJ�J�-��4��G ���RJO��-	�`t�L���X���'�G��ŗf����Ws����S�t�@� ��E��
�|l�Bx#n�r� �{�sO5�=C ���'�KQd!�����b�J�0a�s[������5�mv�M{,����k���h�L�in��X�Xxĭ���ì{��p�Ƹʃ�e��e!S���!��"��������VV��`����"70�}���CgX��
W�����fƁo�ZRB{�bO�S��~b�ŧ`�8�`�A�:Zq���,m�߲ŷ8!w��F�dM��S�G�d����[��3���Yz�Oj�͍":7��o���]�O���+1�J��f���SS9 9@�|^M� .�vj�t�`i��5�A����ӣ�8_bQ+���]���V`�gh�
Q�y��ή+�h�|��y,�2��+ >�\�gἭ�r���ul{�ۉ����_�\�1�A��CѶ���?����݇E�T[s�_)S�z��8��Bf�[O~���B�n������D<�D�r��h�,�^�)J�O��O��w'̦Ñ�3s��p�o��=N�
�ov�/�&>�T1aP_|Z�L𯱐�, \�B�n$�Κ�.D[�yYl'��R��M�F%�=, 9A&"ڮ����p-���c�߻�Xg\�۰Y�ùv�ƞVܻ�rZ	s<�$�4�)��7Q��dy]��c&Uǁ��/��FF9QZ��(r1S$)�|��hGO(uQ�-C��V��m��X�:~"��J�&��ʥ�)@����������9ߘƾ�S�2L���W���?th�c�8Ǧ\ŔB����" ��Č�bޙ~�������T�37]�)�W3/�~Cl�0����.[Ю�)ǎ�k!ꠎ����)�U�$���8]XlI>�N��-Eё���h��Z1 �����>x�8�˺�ܶ��P��#U�"y(��V����Y��I��Pj&�2�K��z��l�4��Y�|��	pDہ«��ʣ5����.x(S��!��h��3�)�#��p)������/�0;$�K�KP�0maZ������Zifu'FW�*���<���"w�i?��OH
��ɋ�
�L�"�S����_V�8�F�)�0tM1�Xu��	=ˍ}mQi/P�b��>M�:��#8���8zϔ6�o=PS4�;��ҴO��<ީ�;������jW°3tPx��u����e��4�$X~�Cg�!^"����Jg��M x��b�п8��c1�{�s�!�;S-��B�����0�Ol9V�X�]�W�x-2ȵ��-�buEz���E���vAhŷ�IsǍ��$��P��S�iY�O����0M��v���$X��u��`��LQ+c�
�jg�+��a�4�ݍP{��u��hn]�sΜ�4�>�G��]�5k�գ�95(B��
���[8�sd����^�+sk��1��Fn���^�y!�7��[b^�PV�OuK��B���~�@ !�`�7AD\�c�s/icKl��͓?k�H���NP}O><HSv;�L	2�QkN6�t��PO*+/��Uh�#a�R�	8
\A��)3�}�q�ᄉTz�L�ISBv|��C�K�Jރ�5����Q��+�c�$I!�+����e��@��9��C�����c��p�j�~CJ�%L�1��7\ň�(�	x@ڗ�J.���=�qL�t�@4����3jTowc5Z7sN��W���Y�.�XA ��dsk�i�=$GL�����EG�j�90�ʣ������e8�Va�k��;^8�jc��i���:���!ǈ,`�Ǳ�{j�.X5M��D�pCP�AF���9�T�k'��0��9��[C	�G��e��H��粨�tҍ��ʢ
��:+8�#�1t�n�	[���W��7~�{r̍���y�>�L�]J��Ⱥ�P��bj��!��S+
����
��j�^��[>hA��$)n)���TI��CY�I-��%�����n咸L��� inF��@,�&�O5	�}��_/� �O��s� �jp1:�!�g��oΑ��5)�|1!}�0�"Tǹe��H��d�H7�zfx.~�QE�y��#��#(�k�<%�p�?$G_���4;�4G�5�sf�ߪ�kXR�u��W�R�d*��8�� M�0�o,�w���U�=�z�܊W�����_��PY�5@w���jo��_����k��d��s�6SC�)U�t��w�����9��-������^Nʸ��'k��1�`�24oD���z���rߎ3���"��'��^��f =��4��4���C���T�?��>K�x6��~����,���GQu�������Ӥ��]z�b�(UB�E���%sS� y������A蒪�r�y2�N�I[=[25�����p�z�h52��}�W6A�!,9#�r��Cu3��#��[W�jΡ���IX���ɚy�7����?Y��9/ёsL�L�]]t���(C���w���O�҃���pl{�����7$����a:�ec����5�}��r�LH��>Ϭ5��*Z`(Y�fw�yZ���Nz'x��X��].��C`N�S�p.���eX.:傲��uL�R�$8�6kF��}��M���x�K?7���"9�M�Ŧd�a�1ˬ\���Z�vΟ*MCV�rF5�*�jhx6�}O�{�C��B#a݈m!��g��,�mTpミ	��z��� M�/>� ��� �_�mJ�I&��S��l �Xs�'<�|�)xf����>���3���qc*�e�}!��s�+�d���C�*2�`M���M�J��ɴu8�k�F���ti���$����4����{�5BbXZ�����u"n[�On��GK���G�^C�)@Jr���(BW�F�k�5�P$��ݛ�����#�G�'}����<_��z����'��������j3㒃i�`��)��~_0���ӦbK���k��4����L_�������(��<W2�!2S���@�,�ݿ���
�x�c�S�Z�T�p0#xE���B�c�g6�H3��p[����qC�"����xh���z~I������.��S��vt�;�B�n1p��d�o�uL���8o��ͦ�ފg_S�)XAm��F�oݑ��ĵ��YʔQK0!<Q���v�8�ب�0����$J�����	V��U�_�\}�]���}f����BF�_�Ex��p0��m�x̔Z����.k�5���N��1ܞ�tN���B7�︣�E�� U��A:� Iekk[�{U��5pAM�7_�l$���pЭ�7�F��a[�����>����� V��V�7��B����`F�������� ƜH�2�� Oب�_��� 6�5Z��$ʲ�Tշ"	�bᡐQ���8���8��JpTw �&5��u��r<U��GG�.�uℝ�U�A�-r����K�c�?R4q����M� 6f	�<���q���L��ל�;�����~������,?o�n~^����i��D�������,���4Va�������J=��Y��A�U$�8�-�[�:�	�ת�l�d����
%�M-\/�"ſl���L����&*7]!���[5�J62�/�"��r�L���j����@��U�Kٟa���hZx��-V�"�Z��r���GdM�D9�K��3f�*��8q�T�E~�	CJbVO���'t65x 
�ɾ�c�SS	`�Y�V�1-27�	{o��cj�	�x��Ձ�<$�$��w��0O���{��5ޗ6�z\�(�R�I {i<R�v�W^jx�S\Ȥ�����ZIY�?���g�����<'*��nw*6�.�	_�����s	<�A,��i���r������,(J����z��2�Kɕ|���%=�FI��A��<�h+��pHr���r��y���#�r��}�앋_�Χ-�z\Ο�l��׆'&.��b�1 �a�O�O��[����L�o[��J�[ Xh6b_?Ͱ=�R�SE��ރ ��x�'��r8ݢ����_y�bM�����tl�f�l-��Pџ��:�t=�B��;����ZݠEt��	�'�צ��C7�2(g��?4t�� F���,U *��xp��=�l	���~␊ʼOf��������-ʠ��᝴��PU�:��O����!����'������?Ll�Kouv����c�"C����N�2F�`�v��)��vB��5���|� �?���_��
��rݻ/��C�SY���W\�������G�����XbJ-y�˖?7���2I��S��XlxVHYEB    4f62     b50/�Y?��������t��]L�N"�yD�}:��U��G@�o���.�����C1=���5�� ��֝80�/����սF��Y!q����
E�VLJ��=�v�W��T�-��$�3	��G�7���ACʝp��kY����^!d �U�*Z5�W��/�zÃ�,�Ə���dw�%��膋*��M���Z�Xdj	��#>����,_�N��� `��N�,�H����Y�j�:����2zo �깰�=�A�����*%��,VM����.���J*�<�%�F|���C��ng�J�&f���y��t$�+��It4}RE!���'x�.S#ݮL�ȗ]+�r~��.Ƭqf{8�):��rL�tK��7!��`7`C�HE�/߂:�+��_��~�h�c�S�t�jb���W8�����AM���+����7�\�s�'�J*�7'�<Q!8$F�-|�Vf��2��2ܼ������ɝ��g�#j"���^f�$pI���y委��X��C�Ȩ0�/����<bUyECIX^�K��S@�\ Cc�Z x��R!*��г��N�'�	4C8�]�`�W���~��|��ՠ�2�d�S5�+�#~�W@u�Qsh9��@��g�����`��Dlʱ���^���O��N����rq=tLii6���ˇ{|¹Yt/��1cDt���O�7Ŀފ�0\�㰕f\h^�
$���Y�c�8MU��:��L>4��}Ӻ*�����-��qD3kh�.mE�ܡQW���[9Zx��!į�KL�Q�!_vL�|�0JUD^��[���{�����S�s�WCEW=����L@�5VW���܊�L������b ��<9&w�M��T^21�g(_"�� W�.����xD��>��Gb(��	*��}���3k�i�B��M��D�q�q�u6�OG�GKwJ�^���N[�l��D���b��	���{y�Yb��i��c��.	��2��5��d��fܘ�^	��n\5;G�Zg=�I6s�6�##�F�qe�E9g�Qb�s��S��R~�o"��u�����Zӳ����{V��p}����U��co��]����V��c\���pB釰[8���Ԟ����v3���bJ9o|<=.N�Kq_&�o��f@�j��� 
�����h5�+�<��8��:�%P�E�Q�Ϧy;rur��|Hc$}��;Ͷ��!Nv���b@�J@o�\7��b�=m�������a�i���?!�W7�[12���m�1,��ZLgx��R�=������=�59y�o�hl�N����L`m�K\��DQ��Az�)hGP��Z���ˋG��U:����|�t�G"�K[i��m\~M��O��[�*�e���g@����P*���pha�E�C\��kb�I�nSH��#�fʲc�vҏ��ZP��~�x��o���H�,\`)A���ȿ$�nE�<�{����ey�>:O���)fU+��??��[
�|-�/�,AАd�'�^�ծ����ݾ�O'��`%Z۸��[�,J���ۑ�!q+N�s�4�xЀV7,�󔬂�_Q7"
ƀ$�{���9���n ޅ�-�b���+�V9���D^��+�C��g���N�B�"�GVP��B�h�R�D�1������7�R����T��'��퀐��+��&:����8%�����)p��$��5au�[ۊ\��N�i^E�oT��8�P٫��#�S	��%[�
�Fiq:��*������ X��%��ݭ�-�ioD��p�_��,�'d����p��ԃ�������̉yoth	�"�$����f����UB�������6i߮>�a�*��B��i�_��k�sn�ջ���cj6��;���0��}}�E3���)4`1#@�3U�Y*���G<Y�b��V�p6-]�vr�yR���sqW^�KI�D�4�X�)�"E���k�Roy�+�<ca����٢�%�����^��܆I2#rEn����̟�G&��b,���ʛ�q��ZYS:7ˡ4'��-��a�o�}d1�D�2�Q*2	M�@N@f$F�A_��p�d+�����<R�̞���eZ�&�v��\;�Lx�,ZR-�t���f���g�l�41og'�Q[*����{�C��\�".'�D\d2��o��v��tـ��e��2G4��fg$����?��\��ϖ�m}*�`q`'ϩ ������X�
�F��ՕwYJעR����Ȁ���2��8�n�?E:����v4�|^d.�N9�?,&'���Ȼ?�(�ጴ#������>����@gŲ�9b�TO	��-�'����50�D���N�X�=C�7}-dԓ����:}u�m&z�4m�C�Y��@f��F��BL����g޶�g�)�5�n��K9Fr|����������#ytW�r��O��%3�^ ٵ�4.v�t].�v�AH�K_�{��<��oUJ�ʐ��Z�;L����R�����w!r�1�%��zϏN�D�se�k������b�Y��̑�J۞2�u���P�۬�Yr�Eň�­�_�9u ��r�q��@,��u]���c�] ��'Y�}��?� ��3�UP�sD�i�jF����x�tG�.Tﴍ�����wh�v�2�MO���44�HSs���!c>6�;�K���P������]!��r�%��r�)�)�7��v3�k�,!h��"Su�t���MǕXJ��R�M��b�9�kDe��P�w�J�\e�ܭ��G�}˅���}�?�V���M�۟��2b`d�D���E��r�B[d�RM� U�^3��Oj�2G�{/.s�/{hR