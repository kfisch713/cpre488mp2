XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���W_s�a��Ο����f6�B��2	���r�����"�,h�9�BM�_)]L����%ᙸ�by���R�!�7[��ic��i�F��}	M����Ugw�ډ=�gڳn�|�6.�\�.D�$sg�9	�Ǣ��Ri��f%?�P�ߤB���O��yu��#��ԷI�f��z{Z����b��y%�IJNH�ur�;�2�� @�3G����b�弇�E��L&!U�i}���L�.�:�@q�8���9�}L(��
9z���df�ˇҧ�����=a\G�:a4�i��1�B�����$��IX�g�sAJf��3�rx7~��C���Z@�m���e�p}�r�ׯ�U3���{�Ri5k}+R,�4��I=/�(Ǹ{�M���W�M��L[S7��Ԭ�#��;�^���Fp|m�Y	P�tX��ǒ\�L3RÎ z���H_Fr��}�i8r������UN�y�=_Ćm���魰��O�_�!J!��w>�Yz�엘=�A�B�+�|⚀RhP"D�h�[�eR���5ɥ�b��Ԭ]�c���������.A���Cl�CH�)��{Ԯ�oN.�_�e�c��-f�f[w�{��������/r;[RT`�Au6e��i2D��Pu���Ug�t��|��a��9�B���b䧽L�F�B�t�PRd��FrX?��w�-��QKU��Y��!��R������؅��c��)U��%4�������Q?��Ҡ�di�E-����)Q�^i�ŻXlxVHYEB    4b9c    1300�:���U��L�7�-��\�ԚCxraR�<p�`�����!�M	��.H��w�B@&�}�q���Ң*o���Z�����A��*Ԋ�Q梥	���'BeV��~ �Q-C��ڣa����s��}A���V����S��h���\,�� P��w��yՓ��K�ɸ�'�&l��Q
=p�C�������ؔ[��q�|"O��hǂu�Op����)Te�Į�εey����P��� k�Mn��"��tM��>�~��~�=�j�W[��"���a���R,8�����Ӊ��A��c���l�Y楐q��mY$׃+*�d{I���>7Z�y��4�i��9�jCɰ��σf��װ�	�QJT5�È�:�.=z<pV�
��vR�J��K'��3��H\@���N����o��'��2�6a���:"������]ѳ(|�w�eY��Ɠ�����!��7�
L�z��4����$�2M�d�I�F�	t3qm��yt��[IV��i�X�C��O��
8�+���B��a�.��\7�t��� Ip�ġ$�.tMւ�^�D��+��	��������N��B@�C9�]�~/;�NH�R,dX��,S�Şc�߄WsX���vҬ�Ar����b�5�	�;7�1~Ti�j�=�~uK��t��>�I����+�n��OMA,�hB�p�}�:��կ-�3���ԗst�~^sK�UȊ
R]���GknL�_�-�5�T���Xm'��������+���:��"�������MƩ9O�o�#�rɞV��dz��J��H���L��1x�ι|D
�1�[[�����j����!��T���]l6���.H]�N!
�c�+�N5PV�gɠ$)�sݓ��:�.�jƭ@+�:�U���IB�%K����ɬ�⦧	2霟�����*!~�A��!\(8� &�d�/�Y��j�H�$TA	������� Mͩa7�c����<���U�W�w��]�-� R��,E_���<�{�T� ���z'F:���:�F�r	�I��2���G�e@T�&����������h|�=z7j���@�2PD�KX��[�s�s<��q���+������'�Q������P�~O6������n1^��2S�Im5?��ƿ���ł�>6k�?��~q v�ܢ��ӫ�:��\~�%)�����^ogC���*���ƃ�/e/�/�b�`+�WFA? `��-������3�|Zف�`�������?`O�0���ԛ$;DQ�F��Z���ɂ}Mx��KirM~FaGF�U]	��s�J�4��l���d�9�g�n�DnR�}��/��Z��B�������C�]/,C�/��-�Q�c��#|3���D��r[J�Mb7Sd3�
-f]P��{-R��\=�벎@�g�(Xx�{������+bɷ�Kq��jq) *Es����X�>�7J}�h�XΊE�W����v ����v�;3�a���i=CVt��K��),p`p2L)8�§cf�ٖw�$M%�,��ٺ�g�i�n��;��;��#Ia����*��@i�a:��"�sM�[5
��:v��USEUO�@@�emr8H��+����f��t���å}y�w�C��W���Teɦ��q�Ä�dfȂ�7�a��Pg�.�O�pQ���R+	�h���A��k&|���B��>�������mT�b\�zד��O���SA������KT�����40�X���m�tD�W�D����X5-����2��G�;���\�`1��(��ŅF����ɷ�+�1��!gp;�ۄ�j�Q�����qq�b�w��[�7bW��B��Y��v����5�1�WPygַT1��⋻��}#d5&p�?�<��o>�Q���8�1�I8�ǘ#Fqm��Ь�"��զ���i�dG�4����P�B�ρ.���[6l=w��^��X82��+s�?hm�Ǘ����,o�;�0w&@V� �$�Mh���U�%��eY�U7���=i��q0�l
� Ľ��Mׯy8̯eR���-���v"��X���M����&��:~�,+C��ǀSJS
+�����Ͳ�TX��?२x��dpd�.��c󏰨�d�zd���-�����B��9}�~�iM�1���w<����[L���&#R�_�_D�w���f�;Չ*尿<d��Ñ:�.m�W�{(�B��=<꒯K�rN�3?x���t�^�a]��l)JW2&�=ʓ���w��o˙�E8��
;Xqcb��y+��0r��]�/_�s�}^m��#��ĽO��X)9W�CK���/�Ȕ"7����n�S�P�4������Z�9�ܦt�
ܽ�q��wJ>��X����*� ��~Wďڀ��]�3�3�T�)C�y)�Ʋc��=�-��M�SX��#�Xǡ�'��#�>9b�A�����ړ�����P�q&�EU.g��͢2�b�w�ԁl�^�N�L��L="��Oh%�f���&��f^�����;��aY���qI�r�q��=4b��`ő�'�	����Q�TP�*�-?1�j���@͋S+��������!Uj����WܓN��<�U�U|A��p� l<�����i��i9�`�;p��C�����@�[�&��ˍ싢hH!h��T���Z��3�ތ��$ٽ�~;Ew� �>�X&���t�/\�g�;7i:FY�E.�d�z�{�Kk��w&���v\_>�<�ƉT��4��M��*�׷m�_��f�8=���������u����0���+g���+0�~0��m�>�$L�8ʇ�
�ҥL��"3N*�3���؁�F4K�t�� q$�!6� *�1G]����ȇ<Jq�u`���\z��Fc�j�4�M�]5(>!۞��0��Lߖ� �����x
7B1�7�>zط���(F�*u��q�(Y��I�K��9�˨��e����=Ь�w���q/?���{��{*��3��b�_a/P�x�{��R.��Vי�p�I�v�.�����ML�(�7�ƞ�G��SBlt��|������|�~@�ew屛�"���I�rRÆ�"w��c�����r�Ҙ�ߏ'8��2�r$�By*�%�itaŷ����4o�61�g�I̟��)�z��f=���ڗ�P�kst v���LpZD\����Uu�����a�j2n��؂�KS�?c����/P��hb���s�)l�Vڗ?���_c&��mh�&�"��!���e�g~&5�.8�bܗ����q�A��x� ח�|��	<%��#[n��:70����DŖ_f��^6�����Z�)ޝb��%�Pn���3'���ި��S�f���U;�� �,��"�k8�'��9����;�"*�d�����>�A�k2Xڌ�u�f���C-Ӟ�ӟ��{ϒ^FE �-�t�������
E�^k���ظ&q&s���5?1�z�[O���UX'>�e��S�˭�$<���p�o�HrI�F�'�k��	��Fr@_t�)m�@׮����� ) �a�ls�:*v.�<}6�5d^�ߑ̣���qW8LHl�=�i��"�	!ik'ܼ{�m���d�_�T���c�
�$*Qd������ 
��G�s~4z�0��x��+Q?�����V�O�j,cq�ŗ5-����~�M�/���R�Z��kxϻ*��T�L��)=�m���V�~�6E�zX�8���Q $,&�	N/uƋJ9�b+֋j*�F�E�,�t��Z�m�F�
�Dzˡ�*�[~
��
��qig�#���H�9}e#Ӗ��0�|iul��)ՆH��%j_c��2�����"�i�x��Nn/�XO�ݞ.��jaL?��}.�=^�D�GJ��R�Yr��V`Y���%��Xx�mA��re#D�혎i=]��~?��oD�GFӽ���Z��4'����_�W�4���a0	�� U�؆%?p\�WUVUĭ 	V�A}�l��e�b�E��	
��4-�E�n�倚L�I'�(iIG�Q��џ�'׺�?���o���e5��h5�P�w�rՂ�:uN�&%%�/�kX��?��^��A)sY�Fx��@2�{=���qs�1g�~��
�(�x�J�LP9OM3�/��l"Oq�� CM�6e�݌ܻ��N�mR2�>;»�7i�2��x����϶���a�ԯ{�6�sup�$������p�ez�2V������Y�/�����,�$�uu�v�L��u� �P��[�[�}FQ5"�YUz��,�4���W���ǧ`�i�z��	��=	��Htw�������፭���E�j�#1�Wm�Y�H�����"l ]�+�_����A�i�l}7|v_�����b��h��o��e���AR?�D`D��� i�y6��/>�|��J�R��FLt�m;�O� �2S��r����F;Y�X]d~���x������V%��;��u-�KkI�`Μ������Q��&�/�$��;;��Х6Yͤ��m����PY��Վ��q�gx����$oC�[\v��h����+��A ��7a_h�>O�=�o�#Az͍�����v0u���2#�G��ޑ�y6�o�L�}�^����x��\��)�b�.�7Id,�&X\�d�A��<�����~?��eepx�[���v5���a�~��oĝ��L[{�|��ʉ����~����:�M�������W!�q˖
Z��v����w��]�e�aUa�`�#��T�{�L���-�m3���8���R%�M��},���/O�<