XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���孴=Xr,�4����jӏo��&"NίO�;�l�k� �`A`�ްv�B�v�"_uݖ��c���c��NX�,����0��dTbUeww�
�G����/���r�JLt����HgW�u+�2����pnO�T^9����_��Q�	�$1��|���/�`����9
i��I�����Th��u��S\�B:jm��d��2�����m�X�_f�'�{�+k�JF����l�<a9ǆ�)�/E��*�b<�0����:f-���[�uhxp�&��.{����v�'C�8���7˘�E1d��h��/j_��b��0��*�!�6�5&fTW��En�C�~��f�bon�Vi��<=�:���< �3K�:�X�W�c�^6����ʯ6K~�V(Y�%�"�ڭn<��GS���d�x/�X�D�Z	�&(��d��UAn��!��
�o�"��'k��XIq���~������2�Oė�!Q��lP�5v��Ҡ�<��pC�B}�I���ɱ�I�l�m�x.�"-y����<0�C�a�P���x�Lt�z:�~��q���U������l�A�~b��?.��f���β����SoO�1��h��!��>�5M�I�i�9H8�������r��;��ph�Q�g!��D+F���:�+5t�`�3ݶA�}�o����{~]ؑO�
��usm�CM���5$�iy�1@_?�6"��:r��mQ�u {�N��N����J��+B�� '3AvGђf���Q�$XlxVHYEB    3e93    10b0�N�-!���~z�5��V�HO�T�����JUX���������i�AoQ���s4�����w(w4XI��o��x&�%��F��&�rQ��\�sq$}�A��2�-S�)y<���P�.��L��P���ǩf�ә����+4���*�ZPm#�]S����)K�'��J�[�b�:Ա'u=�B	�A��1�uS���s��22Y�G8���,E:n=Qߣ���
Έ+�?�#�뾆n��>�!�8�����/t�<A�.D�$���:a����b�)�ZS1��|p���nR�-�g=yasU��~D�����h�m�B�� ����#����c,I��ʊ䳌���?��X������~$ʂ+�jU&R�t�\��"�v/������Ј	Tv5p�����_*LHI��͘ޚs/v��6�Q÷X�({1��)���L�2_�y��:s�r:�����Put��K����ql��(��9�Ku0�\�zח�R͍��#�3����"zf0}D�wZ�>�W��ځ��)���+���e�E�x����MR��㤣J�Ϗs��'�( 3,q:�P@H��^�ħ���)��a�Y��R��%݀�]� �hL���˽0i��U�k��X��"��#�4�<���"#A��Ђ�o;Ǩ�U�2B��'�e�ٯ���S]��)��?O?`9�.a���o�8^����G�����	����ӧn�Bg��i��)r�u��nG������)���|� Z	�V���5�1,��d֤d�j,����v�d�BBU�p�G�B�g���-;fQ�u�]�*"�pO��g$$l(ʷ�K���A�e ry�mރ���-�of�=�P`8��|����%k��P�12���&Ie�'�$�P������r����K)e���u����F0t�v�����UV��2��,9�U�T�\�5a�jq�Dx۵aL�����Dep:�|����FJ�iM31D�.ȅtА5|�0o��L`f����(g�ew#s�ힵ�R� �۟�\W�7����t@����8���A��E������=b\t2��,�R��ðk��g�f�?>ү�u09�:�T�V#����h�,у������R~u��ּ�>����~��A]_�����?�Ձ��~��ǜI�		���#71t�7A��,��)ZP�t�/�ɽ�ɕ�V� p7����-����*�K%�V��mw׮K�!�TՊ�Q�ٱ�WI�6r�U��Ww���+/�`��|���Y�u!�6�
b���cO�_��[�[$y���]L�8�*�^y�c�,��)���������I�]�Й#�][\̩���Qf�Ubҵ�{	�rWݗe�ܮԒhD�����<��� ,�F�Xq��z���A#l��6�͂)#�Q�E�Ah��$�z:�A��/�S3]�zA/Hb�r�>O��������_���YR�`�U�_���lӍj"�;h`7L�!3�L���p�gϠ�c��M���4q�c�!��u���)n�y�������D�n>�6�_?~L\���ge�6��/����B��3U�l�fk��z��}�
��c7�|(���˷E�y5Vlޥ�ꮲޔEe����J�4�+4���:�PW[�ۇ���	�%�9���p;k�镳�y�7�z��s��=
�~ށ�<����R�3３���.��:լ~�>��t�[�q�<�+��Hm^�S2r�,>~kM`�`b.�z8�MpY��P	��f:w/ϭ
���^�L�A�"C��͝�P�d�/��eS.6�q3r�nmm�<Б�	��ᚄ�t`1�C9��d�P���t�W���?�}�LM���#�¹�blw�Sl�D����D�$���4m��IM?*�<���9�\/] al��b�|�'=:7�K��ic�§ǉw��K�c��7�?w,3��ަ��v�9;(�ݞ��N����E�����^�H�N>���i}ߋ@���ey�fu� ��h�I뎞�`gm"Lz~~�y�6�~mr�y����ư�N��vY0�J���ʊ.�_#K�N,l��H�e(�r��B>�Jyw��u�B�BSz��{�^�3���<z�.%�+&��R��)�&���`�Dp��`���ŏ�
U˕ɍt��32�|��~�����,b��� ��y"�Ԭ)��1
�Sx��*���Nb�@ԏQ[�˶�	 �����[VQ:�U���®�f�]]yV4]=v�Ciu6H)�,�/�Q�����C]��ioƍyl���'hI�;�B5�+=F�dg���W�\��Ker����E��/��),*7q����f>��h/1y$KpL"��P�X��eE'�S�wJ��&�9�Z�A]x$�-��<���2�1@u@�x7��ShV����^�':,~����_�.��"��Z���bq�g�uC�`��mg��6��mn�K�i{���~��[�9���܃��W�;�%*N�C���Y�7�>!�K]x�σR��XLpą,"�H�va"�	�1|����8˳�����v`B��XcH��Qq�J�M��>N��Ժp{%�0*͎�ی�hC�\�BϷ��E5v���`�n��H!��%�SHHA��էȱ"�z[P3��j�D3(l��!�����O[f^�E#\�����{#}��q*V��UWs�R�7�ZQ�މLB���h�����<*Ђ���U;�IeCÞ;�,A��6�Y���E��o<�4�^���yQ1/���<:�ff@݉.h*6{�r��h��Ŵj���kv����=��ů$#v��X+Z����*�#���9�$2�>?�#uR�U�N���r~+S5C�,�ˠ���l�Zo����2��{��*��!b��W{���stm1SƧ�e��-��� w�'�u���m_���7�����1y65:�)1�L��Jz�N\�a]~k����l�Y�V�ؾ��j���������L]z��`iu���s)11�(� T�9��&1�jn\��B�ST���^)�)��s,N����ӌ���oh_���B{[�Ntj����I�Zl�,܍B"J����J���ٞv_S�gA�\L��[(�t���Q*����P~!�N�G'[�b?խ��B����X,�r�"s��^"e����戼xER�F "�R��R�f�=m�'1�Sj�$r��C}��R��0�w�%�p0��2ge-�q��O�m�f�~�n�I��q����]t���D����ز�ʃջ�\݀�ڬ!�S.ګ(��V�G�y�A���6#U�,x��}�/dkE���Y�������vW6������`^��Vd|��<��e˲�
���+o�E��p�0՗�zt�X����׏- ;��.�W�@����j+�M�`"N'�^�E�5H��K�i�0��H.�ɛݎNI��9P�dF��xu+����t�D1�!��֓4�W��1���<!���z����Bϡ�Ox)�Tl��i8F��(<>'H�3|���<95b']N��ᒕ��y&��b*�b�b@CV@̿s�j-F�{��y��[	�����ئ���ji{�.�⛗V+�u���j���������uG� %�T�Zb��9w������D/&��*S�U��Ǝ�M)���i���H_'pC�>.����W���m����(�2�Mjp�o��n���d�����e�/VP !�`���^60�BCy��G��Q�&�d0m߃�I�Y�3#A疙�	"�3�19���8��(�(ݜ����4*_մaU�Y/
���2���~ʛ�R�]d�-��~�fǤ�X��br("3���H�_Ǵ%cB� \;�����+hy�9⾞��5��P1��;tw�biX]�5¹~����m��E��4����ю��5
l,?d����RX_d�'�$��Wв��6֤�s>��cԈ��/�.#}"�ݢW;/ 8��XO�����o����$�:5jI�أN[Z@��BD������Xqȉ� �U ��=e�002�v,b7��|����
X+��̼��i#��^�r� 4��ꃲ���wA6.%C/���3<�p�kr��dW��1?�?�F�ZĚ�:p�I2�Hc$[���O��g�R${q��
Q��<������Q�0��북sh����14
1��w����~���W��?���g�A����s�}_�Yϴ?�!��觱ߟ���徰�y�/� 