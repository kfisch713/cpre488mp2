XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`?W]��dSK�ǎ O%�Ipd�`�ὀ��7��|\�L�Ys��gw�\՘�C�%��m�`UN�亠M#��rO�:YsO�*y\/�����ގWN�"�����V=B���=fvV��eO[]b���Q�*ƣ��S�ڟ���U�v�yO�\��͐w�������.�������S�J�O�����/�g�$�ɴpP�B�V�EQ�H�Yt��,G,��u��ؽ�b�@�9��2�q0T?��<|X5w᳹U�Ӧ����W��� ��#0w
��F�	�5�=3��ܬ��|'�jx�	�M	X�0rC]sc�-l)�Ȭ�Ͱ�M�w)��� ��ԋ�w
�nNxo�2�Z�ܑ�jp�����s��6����:��	M�؀��A\�J���
5\�d�K����UY��Q�ve���UzZ����	�@��q��TJP̄O& Q�R���Ly��mBE(E��������=�́*�+�����T���+m�ᱡ��Ω�ᛡ� ����|��l���C�>ly��{~5!%>��Ã:m
����a� #ԇ�ʮ�H��6��cE�]�;�y��+fݤ"[0W�F�4�,,�p��0�~3��crnL¶���1}��2��HfJ��M��+#����t-O��~��\{|��М=��o�y�K��w����8����h�Vm�� ��c�)��1M6��C��_]�L�׭�s�ޥ��Xr�8�qU0-����������Q�Y>��Wo��C�
��̩{���XlxVHYEB    4052    10f0�\'�EN<��S�m�2���s����U�S�mTm�����(�~�V�5;=�wΘ}a�Um��l��LCU�Sn	�3��-E�T��;҉��}�#��?s��B#�{3�"m�-�[��C�� B�n�.�����ɁK�O����1Iˤ��ᵧ��O�P��	U��}+Hq�4_���;�?��Wz���F�Gx	�)[���S+�[[�7����lR2�9z!��6.��FQwf���:h\w?:�ie�6��*)��~�L?e!�ps}���);kA��?o���q�X�/��"�ꂑ�I�$����]ϘdJ��B���+�Y�`��p�t����˂�G�5�Ϟ�&Na�v���ڽpŗ��%�����@@���t���"���5�t�WO��b��҇}e�^���<mjr�R�[����ܫ�6�9��@�L���Fc���Hm��N]�q:*�$\7m
��r� R�������+������=��6\nb��O����z-+�J �p*P�# )P=��>���N<�Ǚ��mF�9�%/gv�
�d^���g3	�-;��#�(#9
r]`�W%jړJ
�6�D�xzW�4�vm�ڥ������ސ�Xm�d��Q���_��	��M����fkP���Ǵu��넀.�Tz֍��u�Wyns���:���q�OoL��<>^40��{��߯!_i�.�q~(��zp��ty̛�l��-�ak�����*yoHG�?�d_����Y���]��,��( ��쐨 ��3�����4�@}��"�DvO30�ڗ�ۈщ-�(|��v�� J�0��߷���Hbt�(~�6�|���M��3+�!�Uy����9D���h���v���~�:wƕ��չ0��4�k�9qj������
T5�l��|��Rl�0t�"��T�剌N|�gN�C�A``K�=��@+�0Me�׍���������L��_��%MIL�-��B_:䉿<�ν����B�s9?N~�%�9�ɲ=��"���u6۠���U�Ԛ�͏fP#�KZ��?�˼X 'Ta\���A�2�h�n�;~H�sk�q���M�cN� �E4�X����θ ,<��[������]���d����^��'D�Y��%N�Yf�4�%�9�`D�|A��*�Eϧ�r�ʇ��������5�An�Y��/�*b#���EA>�`|��W@�#G�Y���w*,}s߅ )�*'�YT.�rt��Uv����d���x����6�aP��(D���pw�{ȕ����E�����+	M��۞�Z>C�I�����or�����M��K[���<[�p���=Q@�l���g~��W�f
���%z(�!��4_��U'�
h|�o4}n�~XMӏ��a:N*���Z���T�֝�VVxEƧ����|����ZX�þ�'#�װ���'a�;]ڽIt�.q���}�|���7O���4�HXĜ-Ie��K*��"n����{�&O���2��#�b���z�k������l���I��k`$�܀ވȈ��-@��ƐN�7��|ӵ����Me�¶�ݔ;u��F+#ޕ/�on�Yfl�^�@nǫ��o*�n���3�#{�ZD}Z�**��F&ҧz˥��-���{�>/�v����,A~�{���$<�j�p�m���}� C����	y�N�=Ku,�9�HT� ���=����Է�N��|��0����V��i��K����ߘ�W�Y�MtF��'M�UoD�(F#9�+�@_U��P��8�F�����Y4)�!e̡����P�'��gb�4Y�O��m6*O`�9��(
sW�����	n����K���D�j^��|!�#�܍�>-廪q	DP����l,�`��b��=��,b���ƣ%����^�@�f ���w��mx�(..qE��h~R���r����-#�MSHg�TS�P��j8����P��G0�U9��ԩ�v�4�n֢�`d�9������
`�� ���չ�f�k��,��/��D�j.C����!���2d�̅��L�8j"���t�9քU���f06ع���I����<�y!~���l����5k�0!k�
�d�-o�Vn�"���/�G�¥T:�.�'����m����͎n��b ފ�_Z�6��8�p�Us.����^����~�U�V�����+��)F.�*���.(�]��"���ii�������þ�8`GPɿ�pj����B�� ��(Ύq�1�?ZE����l��S�܍k��쿶�I��V*��F8���xH��1�8��99�-�JֈJtw���
�,k�mb*P�� ��j_� z4�_ݲ\yq���>��#9����M=V(suc�[.m�1,�|1aͧ>>z�:b�mB�~���8�c�����w|������y��Em��q�Ӣ���t�S�咩�G=r�����ݦ�����E�fp�g��J�M+9��#��Ȥ0�/�E��< r�_�^���� "���y�8o��W;�B(���.ɜ�S�0�uaȑ�E1�F;���Sf�"���ҴXg�����};-���eה�
�����[�����p��){>���:��4O�aaiڈsR���S�~O�VJO���k�#!k��_�f�<|<�:����
�i�Ȳ�)�籥���6��)�ӛ�{�^"�4
�����H#���l�E\1z)��ȅN)(Ix��H�7���P��Xm߄kXO��Ni�x���8'˙r��t\0̯�K���S����u��LzM@x�M�DZ#�O;�]TF�k�c�At4ƒSM�d����p���i�}��3���c�{Hi��O+�`T[k�oi���M�K��y"l���yx�9��<��+K�h�s���4 �V�$0��X(ea�A����|q�����{�F���W��x�ւ��A��zڭ�w�-��J���U�č�?�x�~�q	>E��T��3�|$�L��7�y
�����1��`�ş��r�$��% ���k�U$���RSD�Pm?UVs��#�Ԑ�I��F1�G�+ �cQ*�1���j�5��/7Q�R��I�f��y���7ۦ�����lb� �Jm:bۍ+@�p3��F�����)hs^��<�]1k��UR(� R�N�[֋�����x�\�\�c�]��-�����L���s��m�A��F/~ϓq��J�0�O_M���Is��045,#o�5k�s>��9��$A���{�tP���nGY����$v$h�S
�n�h"���@Ѣ�	^iY��!t����O��S�Վ���;��.��N�}�\UAB9R���{��a$�g6�<�̔YR4%�=L�9����qY�e�f��!_>�D�c�dx��~>�7~X�f���r��>~�.�0�.=�\�Qxn*Z&��9 �kff�zk����t�A2�Ght��Ե��lv�N4J�Y�����~zG�Ь�W��u2Ĥ���멺��Z}sJΌ�Hv̔��/Zt����Pۣ2���ϥ���~[�G�س	l���b���L������GeZzn��<8���bN5��{��^����i;�{�eL��=��]����I��1[#ǖD�w4x�@���뙟M\�]'r���6�`5TB�k��G���i�E�y���Qކ�Y�0N�8(�Jr�L��i��n�d��Ga�O,t�c4�:���{-�� ��	>�;�L�s���~�Ȧ��%\�6�/3�PI"â�će`��;R �E��(h�k lV��^�Av��;���ys�Q6�I[��&��r�����'k��8�n���{E��G=<�T�����o_��ӭx]�1o�_��t��s�������y�81��E-�4���O������O.pMݱ 2ۇ�[8
�M!)���kRg�+K�i��aiϏ3��G��Ds��ȼ�s��D�_��@��������W�Vof�D�J�cQ�n8E���a}}��'Y:������jyt�ݩO��X�!t��q��$���#s[4a��!����ip���[+�c"�ʉ�V�xf �	��\��;�9��,q�oC�-��_Am_������pLKq�^�TQ&`S���`ē��>����ˠ�-�
�쾛^;�1�p���H��l��@{<�7���[� �k/ʀ��v��
��uү �D7�H�����>��|���� ����X-Rf4�G�UU-:��c���,�n����3N\h����#��Ͻ%�|F