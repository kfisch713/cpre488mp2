XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0#���р����cȖl�6��ǽͅ���	N�RQ�`�驕*�㎗�x*�{�����\f�ׄ��_!��5�A�㇗�Dʙ�,�(׀�9�T��B�<9�����8GI{���]� 6�+�դ�)v!ڟ�����W�o?۝���wP�$"8�i ��^D�����J-��c@7d7��ló��<3<|�`�q�0-��G��/rj#��}�;�ߗ�`<�x�d�C6C`y?Ֆc�p��^O�r��;솭�f��VP�ak�ۨ��
��ȧ��"9%كOX��쮨f��T��z�h�4����L��=�����o��!�p�Uį5~"]1)A����L�Їb����9��Y�H��/�����]��4Ϭ�j�#�0.���9�w1�2�[��`�G��C jw��K6�s�M!�!�4�E9���KV��]E�8��� ����$;}#*��4�u.��S���!�A�a�Cy������NRpz�C�a@iC���To-�]	�'�-%��%^�(>dW��	I6�۔������!K.*8H���z��G��ՂX�����[�o.���_�oAb��-.ڼJ�"���ѓ�h!V(�"|WM=���q@�p�Tn�٦�"r�5�%k������^!��/���Q�t���E2�G�6�'Ń�Q6P���~��3��4�1 �h��˒�>�lV�RH���H���Q��s9��ιzp�5�E�S�G��+0��*X%n�ڎ���^f�(��.^XlxVHYEB    1448     800t�cѭ79��0r�����B..	&H�\��[[�����:��;@}|���ט���D5���/8:µY�lh}�>!æ0!AH�8���ust�A�b ����6�8^\b����V�69M�X����.�̧Q��hҶ;U�]�9�����q�w�Gz��������3�
\�H�E��4xEB�ɳ�J�ri&���aQ���>���Q�,�
p��X�3��u��r*=�\3x&}§��a|nj	�y���o�sN�:�_{��]}�ݓ����)�1#4�E����E0@o�黦� Da�������-Z������>.�BGN�]&�4�v��x�R��%��㪝Wa�>�������6'\>`��p�{�V/�T"�v��T|TD����\{��#>mlZ/�b�G&�����%+ -avOJ=K��j�r@i]�����+A��c��j_�2�6�����k`�*W���O(}�O>�b*<��5Nc�jȇZg�g]��BCۃyn[\���e�ڗ����D-��FW;G��B�^�w�1�CKE�Pl�W��ZG,�޾Dv ������%i�0{y$���nѰ�<Si7=���(t?�7M0����%�:���M�3>������e�Eȓ}�p�=.��\{��͗�T��u�IL���~[���]���Z������xs��GFC-�Y�q����ԡ��0�V�G���!0��x!��}�֯�c���j���nE*a��������_��D**ܤ�]r���'w"0�����"�_�WI]��&�P�o�����M��)��Ev�ۯ���/�ˍ�y�>���������R]��4��I�����c�����]=JG��!��}��W���w:t�h�&5���?Z����'b;Kͥ-SӢ�}�"R K��'=I+�Z�=,J9�_/�]vU�2��@�s��!	T-�?�#�.��W�R̂SI�A:��cc���
ҏ\Y��g�ئj�uG��׆�ǖ�8�Z���I%'+���w�S��簱o��g�D��?�V���$�z E�-)�ed��j|F��_�X��H8PB�p6O�-��i��/����	3�~W�./�"�eP�'&�	۪�� W8�=����PU��S��2��%xd��_�Xa ������=ӈ�)�\�WB���i�l*8"�Չ�ݚ���o�Ow���]�lFS^%Kh�+��gհ�����Ȣ��L��R���a^�'/�aSO��'KXkg�k���^���G�+��R^�HU���+
o%�'E�M����0:lf۞=W�e�&4es��~�Q�W�w��$�~O�T>?@(�/�dPC.01�Et���ӝ�J�w_�Ea|I�`pD��ߝ�vF���6��j8f�ϩ����Z�U��΋3ժ$�����=8�[���*v�N���G{��}��{�<#�2�f�P��	�J%�~�̵ݙbj ���`ݤ)~�*.�y[�`ǟO��p9��w����{r�y�����afj�"�'���a%FG���#FZ�i��y`���`�2�ʒj���1 ����|�U�����I�3�G�23�d݌�3��D���j�e��z'`R�<d���Cˆ��n�b�U������[��<k2�>/i���
2Шe�����p�plps���x.�  d��4>���t^�y!\<���{���϶7�e�XP�;�Tެ�=ϛWp�{�,��c�����i��~݀�1��V���@8{3��Y-N��C��ް�=��{�/�;o������tB�*��ǡ�!�t+o;��g��7�F<�G�@����cɷ	�hR�/�`<���F���F	�2���;�F�J�z��y�6�ĠB��,�����>��ׄ
x�J�ID�&��/���;�}�>lמ5Q�/Q~� �p���kȉ!M-��_�ˀbN�(�|��&�4���7��ŉ4 7|�y���;�t���4��;�sӳ>T�]���,�G��