XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z���o>�o�����Ȓ;�̶O/�d49�5�yp��D���ϧ���(�$ns�����L�΢��Fk���R}
�"�lI�2G�+�ƍn���3e�7niϝ2Ǣ��`�a����(�Mh��Ñ!��.�J��	92��K�| �9{4�*����m��TuT�t��K\�]�E��93������#����M�,dj�WWO��9�q"���ɹĨ��f�gWS��y�S(B�����gU?���^���7%��M�=W�tқ�䤤��*c?uO��Ta%/ڋ���i��WU(7�:��WEg3 d�ҙ���Ġ�#�sK�ܼ�)h��p��:s`�\���>���Y��OP�l�R�^�����S��AuFN�6 ����'T	@��^��*��Vd�W�|�$��1���#:0IȔ₺�䍳��ÛO���q˯����~�E����v!*��Ƭ��'1���"�1��;�ak��v|/�Ѵ7�8�e��9�MH���>v���} >}�12̇�ta��B�Js�b��mO����)��[��B.��=C�љUf�fJ�ؠ��PYyP��aٙ����@Y�dM��m!�~:��+�|;��WT� �'�`w�l�
��P�]��
�0��A�
�ě�N}�;T�_l�oŜ�h�/SZ��u�y��F���,i3\%�`�Οd��J���5�R��un�j~̜���n�){Z�RB�w:kq����~XlxVHYEB    48e3     e00���KܶL��8@��c����>�2I3�
RR�AJ�&���T�Wp��,�J���,I�"�fˋʏ�P�(��o�;���1 ��=

8�.�����wB�O�臇��|�g��IU�V�瘦h�b�����Ӧ�l�{R��	%�ޞ"���X��*l\�<gK��X�]�p�6a�+��*g��
��6�`y!�Z�/�հ�VB�>*���W���V~��؆���h��T��s&h�%��>�S(%P�Y��kv��"�Τܗ,��5ة�~MG��l��%�G:DG+O+R��'7�����Y�O%��Yӧ��$��m'|&����Ӫ���ɍWZN�̌#WP�F��w�Y�&(4Q�c'�a]l]�#�M�-l��!NVk��\6�	��z+�#Pe��$�P �9���V�����-�dMm�[6�K�����s�o(���%�ۧ>�{� �"B����=�ү|U�L���_.R,yT]`!�E�lZ��%|��Jς6J��^�}{x\��n.��
�����26���`��K�}]��qy��~8:}ئ�����{�`�f�7��F�gف�Co*�!wme��h�;�y�ݳ�)�+��Aw�z[���s����P��������	�;�׬ �ݫ¹�X�L*W��?�D`Ul7�В#��F���ZE�`*xa�d���� ���e>o-��x�^�����#Uj�kR���-+���sw��-��)�3!��d/?�x5e����	�Xh�Jb��Q|f�~���f�h�H�,'����O����H���3uW�>_�3h�;�"GW�
̒A*S�����Vt�,�	�N��xoR7�$���G�c�Wk<|�ȹj1�_�+=�6�^���sP���,��#��mf�w$�h)z�g�����'��%a�P����ڳ�������:v�]�¡�#Y65�^�31n�6��*�I�=��ox��5td�5ի1�2�����wW���w!�o[�W�>��Gu��Kk
�Y��pc��$F��Ł���6�0ڷؾ�)���oi�r �G���M��S�)�=It|tql���8*�e��B�t�ʬ9A��_qQ.����X���5�5iS���h�w�4!�rn�
���6��q�O;ط7zz{6�:�2D/S����D�� K��, �.a1ޖm�Gk$@��7�+��Z�+���k�ۧ7dVM�Zzg���D�8�on���$]�k˘����ݷ���'�c	���"���z�T\�p8�S��#d7Xc��c�UxN'�Y|rN��b�͖`���ɹ��y�PqS�z�d�?�W�8�@����C�`Ʈ�u�s���g?I
��R����5�Įȑu����B�u�@����C|�m��?5�H��*7��*K1C �"+M��Y4�U����OJ�AAs����}?��b�U�ZjuЯ��O�+Yɇ�@�}�,��n��	�o�v/���C	�Ys$ Y����Y덭X��iǚ%�(�5�ˠC�c�J�"ͮ�f�*0*��+�[�Ҭ�!��9���h�<~��8�5)����_�;�����b��QÛЩ���`跤�x�!}�Y����)�S^�F�P����[��,�L5�`��iX򽭋]	N �;K�μ1�]56�f�م�fm���[�|�7�����f��n7��.w���tW<���R��sxt�K��!�x�TL�-�sdm�[�e�%��QШ��ru�������y���銳�� �����{��& U����t[�%�眇���>_�\
����v/?M�b�v	{�pY����Tͪ��H	ۍKo� ����ED�	|P�O�=��T �q3!h�
+�*3	ɉ�W��RX#�����F�d.\���n��_����?U��� ��a<��#j��7���k�2h+h/<U��xA�@�<�]
���Z>DW?���X�d2��_.E'e�+KW�-''�0Ϋuv�7����o5�pVV}����֨Z��z!��n�LpJ ]JXXR1��׻d�B2$� {�Ī��iDU�ű��?���S2%668cY�_>������Ф�{�F��E�{g��
��]i*�dq͵�F��݊(��P+[�]7�	c�&�L�=�*������'Gw�
�M�tptG�ajt��m���esxM1��74��%E�	��2���BU!jH�h�7���q��+iჾt�Uh�\d��	��w՟�B�̿�LA�}dCA���}���v�':��K{��,]1f�H|�L�j�(�r4H����/o$��I�rV�Dg�A#m(�^W�ʣ�������W�&�"���������,^�r��g=����8`�7�1�f�����t�B?F������,`C��@����.�EK��c,y�e����꟨���AO{�!���t�GW2!]�	�����\��)��aS��3{�4/����O�>Z�xM��2�mD�M��mX���F��O��f�8�_|�_CoA:��nXp?l��|���q[!ՆK��}��㥘�6y�JZdy�Խy�֍�P,��ڎ�4�Ve�t9���(�B�<u�m�l��#�:���	_��?!����y곿�O��_��\N���~/V�Ż�J}B�����@)f� ���'ҥ���ȃE]@���D9�H-'��s�����5z�OS 4��ok�����C�S��5��n���k½ �n�t��:�}��=����꽁�|����BL��b�Ĭ�wJ��3G9v�/Px��W<p�_�T��H�x2��?aH���,/"��E㧢*�����e}���y�r�4I�'���mƐiv�R��2+��ж�iA��G��o����+�^
wE�9�Mr�\���y��:U7�qG�������s�}����Iy����߽a�z�w�:���g>����=�A"�d�0��0k�w\4v��gf�b`.A�U�]�oQ�R�r����x�re��a��0}�U?���k�I�T	�w��l!�\8��Z�+	b�B�40�I-���f��>���ݕ�'��d�eM�������*���gG��P�5�iFmֽ&>q:�z���%k���~]�m��OR9��U�Y��p��-�p�m�x�]M=i� 8�3��T�:G�#���k���i��`4�_1�<��]/�E��F�<6�����(U�Xb:�M%��?�D�D"/�B���hI���왨�����H�n�B��%�UNsH�$�ݬ��������m��S�(����{� |:�v�%���]Be�e�c���l%��D��j0r85���FnxL�/�OQ����u�p����X[�*vGX�J�{������dk���fE�횐a�:�$�$#���ѣ%���/�M����C��=p��[��k�H���y�����+ѫ�fҷyK�{eC�s���֠�hjǱ�t�~%����	�;�������c�Ը��`��g�p�Ev�I��X���HP'v��-[-��k��u�Z�$�~b1W.`��(����A�0��E'