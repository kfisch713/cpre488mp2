XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bi�������c9֣:RnMɛ{#Y>ng�~��sM��Y;B�D��4l)�9L�e꺮j���wo��(�o��a2	[�O�D�����ࠋv��[�*� �A�� ˉ,����ҥv.�A���]�1Z�]҉�RALR?�(�?������e�m�F|ݚ�\��@����<�����}��� ���8��$���֐tP�C��-D�&�����\Z���ř¡ z�g4ݢ�@�ѯ?4����+�M�\9��#�j��3���L���ܒ�"���7�����F�NTν���*G�`*~�{�"��p�K�Au��A�d�3MԳ��}ݳ��[b��|=`���X���<���`���)���ţ����h�׮���1h�S#&�R�ҴRR�nT_/o���I/�p0���0A����7����f;=�FI겉�Mk��w�_���`(�a���H��G�Err� C�(3{�UV.���|6_��n{����Q�zğ-k� �j����&	����8�b6��d�8� ��J�o�K�?ZW'�E��9r�r�N�q�W֔��������*1�߾�a���(P�� uAOn٭�X#G'�iĴE*B@��A���{`�-���i�r�@K�X碥�8B}?Nc�s���j�_
4�"������_�O��h�"^y:�D��E�j1�`)Z�=��  ��d�T���$,�z�>c�$k������0B��b�	aD�a�*S"�|?ZDe�6R9��(XlxVHYEB    fa00    2a40��X�;���<.��!��{��bxsIS)y�Z\�+w��Q�"5�J�=q;G:�|�{�y�٠[@S��}���}*1��dX�J�u�W� i.5|qO��h�s�3qS���|��!78����c͛�F��������h��!:c�DBJ���a���b}W&�K��P���/K��x�\'�ӛh���.H?�� �#��|�b:�;\�O1q�4v.�p}j 1H���G��T.'�#�%�>a=^^@���<����2�2��6����l�f;ؘ@6ɣ�-�S�)s#�t�z�K�{M�n8���~���ԭ�h��!���A��1�D�]�7�1P��Np$�Uf�bFla��?!8F_�T��&�<�z�� �Z�ppǛ���|��"4x	�>h������	�  �dv�bgF�5O�"���@z�c5�;�>�;}*�j��������"��I�#�|�5O�V%}�/X22�[p��Lגb��Du���.��9�6��0x�I3+��� ��9��6�ZRE\��k?��7ݿs���,�U�֐D�!�A��_}5��qK]�"5�i������ � �mĶX�و�+���Hp)"U�)땢���M��{ۼ��D��~��-��@
���՚��]޳j��(am�(��ߓ_V+���D���)I�����N��
m����p�:Z=�E��d��"o�ስ�s��~�m��v�b=�k�6�x�}��"�|��]r$��C��/4,����&�j^�]ڢ���K�{$R��S�n/R�c/��)����ڧ��ɛBz�+S"��-v�|\��n�~zSXC��ؤ,(�E�m10��+���/R��G�����oǿ�Ha漌�g��Y�#�����*s�:�K�Ϧ��/��N{��pT�&��.��^vdO�ܔ�U�)WU�ּGH�����V��=�m�P�5d��^v�c�����C�ey=U��\�;*瀓��Ř:r{m(ӝ|��L�u��{�nU�����Ij¥���><=�����G�F�8�9���y3Yɦ�Hx~c!V��.:�ʅ*E���g��n���_��\�����7�h!��"��Q۟A=��}!T�ׇ ,焆͓h��s�+_�Ҩb�0\U�b=b%%CHBtX�%X!o�!6�^D2�]��rğ��s�hP��e�<�����=�,�E�Zᅎ�Q�'�:+��
KI����ط�M,&�{��^_�[��A<�&m��b�g�
����s��+n':�F���㨰*�`�)ɴ-��x%�M'�aiB��<�BX��-�G�(�nmg/�6̺4ZO�����i�Ϗ��Yaл�v�g
i��U��m̰8���/#6q������5���#�`a���]�����p����U������?���m--UF���g���p�f8���ʍ�^�ӹ�� �3G9�W@pԴ�Q7:��\�o������qu�c��/��=��k�SP-�t\��j��S�=<�@
�:<�؏��,��73S|�s����N�C�Y���y�����I��g��M_�l4G<��:@��.������	��)d��f�*%y�F�(�H񢽰%r0��[/"iT�x��Ӌ4�Tj��V�q.MҸ�x̹h(���$�N���,�B��wȨ���+<H@��� Նj ߄��hkmtq%�wg�
2d��&�P x��y��b9��HPJ����?�5G��u(�ٰ�bL�%��p���"�<�}|�����.�(uq$+�0�f�O��_d���C�m�Ȁ��iI����b�^�D40�Q� �K�6V\,$��2�3̝f��3�Y2���R��T��@K|��(p;�(O�K�zxg��GB1ڤv�ҷbf���S��������DjY6�6k�OǊ����5uc�A���s�� 6�Z�pX�8U�epzJ��cP��Ǫ�����/�J��5L�(i�v95[��[^��m���\��9S�!�<\ލ+3{4������;ݮ	���X(u1�[ls�� �>ed�S��{3<�2�;$L*�٫��w h�6YY�r��V��M�-���
c��� �VM�6C9�b`W`%�h��ڊ]v����qP�����u���᠃lQ5���ɜ$,D�л0V��H|�L�U���gѪ�(b3�kޭt!����8A�������W����`�i�; ���V}���{�mk�pD[#���]h۽����i$}O�Y�?4[�X�V����1G;����M}Z�r"�ճ�<`��Y�Ђ���Ǆ��K9i�'������R��@��]����������.T*�0��:�����{!c�Z�2DRVD`& ��Ex7��zCۊ(75\t�i�C�؅]-��$�7E者G�ڕ��[�3�~Ow��J�iR�ŕ��^+�p�q��W���n/�� ��ό9����|!��X�	��)��~�C#�����G`�
�X9|/�>pD�D�\��xL�U�a��=ѡx=�����2įɏ'o�{�rB��#��ͅ��N�#Ҭ��DG�s�V0����u�[�u�����'7X��X/,����F#S� ����Ɔ0�jT|�u�S��tǫyw��I4�,n���~�hB��N#�1J�ÄհI��w7�2gk:h�����#o/��AR�~�u֟�q���FɌr��.��`H+�7�X���[Χ�:F�S���̺E2jo�V`��]Ό�=�\z)TY_���º/yG:f2�0dd�8�Uh�m5I��p(�A�kۜ��w����smw���)���@� ���;&��l�r�j�)�`��kގ$�`\�}e�/|_�'� T7�v�7�k��8�ƒ�^ 1fJ$N\�cq���������.���t�<FJ�}�������\ ߱�y|b􈗃a�5�o�{�3;����<3�	�ԵX㇓>`�.�L[7�t~�*�+6�� �~)-a�c;G�B���K�E�V>_��um�O��OM�֠+��.��	&��扳�x�-���.��#�����V �A'��v�.���qbY�{5��\0{���]��YK��͢�TpJLGH:W%�����.[�6�Lzت󖞲�~��o���!�j\�L�?��ԙ����i�@��J>�N�"q$���?�yꋌa���F�~��bD�YK���7���'G�v�����T/i���Gو?��SA�f�]O��Ȑ���X����JD
��T��9������k��9��%EqU�\����c�M�v����^A�х�q~�w%�1wJ��q���d��G㊥ ׿����ݧ`נ7#Z�u������0z�I\(�H"KQ��1�AQ�
�.��ΰXP{&�;�ϣ(�$�6 ��k��R�FJ��du�"F�Cm�j=b�'!�u��n>!��&,L��0x�zn��-�E�-�ıOI�t<H$(IS�ÂM��@��E��v�*��bJ�;���SH�l3z􇰩�O���s�q' �v	�u�N>��*"��;b��$T��	��[�Fm��loݤ�'<��ٰ�K�z2;nh��:�4D�`�XT����3i��?�S���[Tzx����.���[f�lj���5IH���.e����E�.<�b��sG-j��"�'�y�a}�V��(�s�6˚�Y7?��G(��q�Y`M"�����q��B�6����?�%/�5!	�,��!K
{6�}NVx��Q(��E3�!��8�.����c��<%��Ի~�Ǹ²��֍��ѽ�����s0��Kɼ�r�B�RO�q�;���	.7�J��Iwy����1/�`�'f�E��c,���e]#�;D9s�U��J���������>D	0��4��n�+=0�ҷ~��b�w��JyxX��q�������� 4��-���j�>Q'D�a��%u�	@�A\4ڤ�O��p��.	]v^�
 ��}36��C3Ud��ψD�
g�Դ��8��Ȁ�l_d��,}@�� ִ2�I���j�ůw�N�v�s�����=�@�w� �ۂ�:��ݩ�*�hB�ѣ���=;)�|a�}.+@���݃.\#o�y�n@H���T^�a����xi���w7�:K��f/����D��Rl	�g��-�kea��ԥ��_ID�R`PQ�Hb["ʑųR5/��MT������ѵ�jg����ԕ��D�BV攸L*c�2N)F�W��Q^4�`�Q>)�.�^�ϔ�H��ul�3G��B�a~=��������6F;���\��84�zN �in�'�?���d$#6�#s� &\�����7ǣ���W*����$d�����a��P��fm�Q�c%���KZf@�x��?(~�������k <���R̩i*� ���.u�)D'�2�{K�����Uv�nﱠ��3�B��������*!��ūS��
��˂:�S�{Y"-�Bz8 w�z�ٕh�:2 �zV�%g銇$y+ϙH,Y�%>���hAnn��������Eh���3Ij�(��,o��mB8�j%�b����i�!�뚝 R��.�,~af�DH��bU#4�s�'�n��%��r�lś����X$<������5]�*��� ��e;���P��s��^��
S��	����
@9��k���߅��SU<�o�Yx���2��a)&b�����~v�0�+F��	!�/z���;��u<C��}+i�K�~*�ȉ�r(�Q��ݎ?Vr�w^r�Ik'Oj�#>`��̃��<e�aC���]�k��������T)�Ŗ�D�?{���I@��M<��3(���$����X�?�ޖ��x�7�H����F�OS*<���:��V�x��jp�X�ڃu��m��t��kRǝr�R��Tj̵�G7��B��%:Nl?Vc�6G/l��$ 1�f��yr�24��^��۠Ʈa�-bNU9��,�a�9y�Z�B��������-�-%K�;��U��Ua-��fjD(�h��@Xڵ�J0d�#2[�ZB���{�uUa�T�[X�$p!�Ψߚ�9�n�茞�:F��=mHM`=�Z%}�GOlX�҄�S:�F�n%>h�P&RwzD=�2�3ζ��z�x����s�Ӳ���Z%fS#&�\S
�gp�!l�\����J��7������e��\cK .Tl��a��x�L��Wc�FM5o�T~ ű��A▻_��Pw���$�]Jo
�&���"�t�m3w8��{g�1�?���o.m@�~0{jF���K��f��c�}t�Kl�4jh�§�EG)��К�q��I~s3ܽ��q�����*�NQ�{o��Ot8�^��jM�%^�ĀTJ4���	h<ڙ�z��UN^��@׸Cb�b�ޓS� a��Z�/*��AWe���7֖Z��=ϻ>���/$��B���Ew�p�A��gcM@E�	`8D����}otg������7'Աf���u���"(}�2*{s��MjN��ґK�*��s �:@slu8к����=�QB�,�K9��Sh{�s}�z�#�mO��D�rrS����E�]��uM�<V�ۅȚ������4Xt�R�H)����Q$�����΁��l�z,a��A�X���vj����4T�� �G��y�}D�1��%iB0�O�v>�'O��#��6��Ĭ�05E���;���ִY#�_�$1Z��``�xn��3�(<b$kuG�h���(C�_c�u��������l�t���m����0��4�I]�&��el�B�u�w��w,<�ܼzc������z2��-�p4��	�i��e�>�� W��O#���qo�
H>��Ǆ׵U� ���}\t4^p��1]�P���{Ku�!�t!l���JqZ�9J��T���3��5���C�(tB��_���cYU�S�)fGv>�K�'�>%�|�=f�G�q�K���y�	�cxg��^0�����P/j4�갵Nu�Ml��Ny��/'�;����9��j��������L�B�w\b��=��e��#ˮ������|u�8��j��� ���@��m/;�RȴeVvp��m���O�q��|����P�H]H�4t��C����t�Q`b��3�b8Xg��T�U,Ԧx���\�a���P�`s
���d#��Y�sg�H�1���b�0$Z��WC�F�`=50��0X6��#�]o�����zdy�Lb�%�'&�c_���wj�}R�Y�_�)��סW� ����H��S%ݕ"郑y�Xn,�'�w�ʹ����a�������}�̡�`�lGT��c
FxuR�e���ve��I��l��H �k�3J���[m��I[�h��^��e�=RK(���|�|x��y�U�5�P�����\п��*�)��GI�.�������ϡ���4����v�Mv\�=[��/�>�pū�v���� µ*���-fd�����א�G`�U�+{4�=4\m��rS��j%��LQ�+�WQ�.������6�a!�.χ�9.f2hT�� 3&s/�؞]E�c�����&�������f1����݆4��q��B*C���W����h=��3_({����n�y+n����N%$q�p�,>A��0	���u��Nc�I�zы�-��ƈ�"�nl�F��b���5B���6��X���7���V��B.��}qT
��+v�ʨb��ț�k��&�L��28�\�{�h�����'����&B��9��@cX������߮�A�1bw;{1K��@�*;�4��{/C9�7���������V^�؈��%�� 8{���{�,�����{H��ࢢ�4��q4�]�E9z�x�ޙk�דx�0h��!��'mi݌�k�k]�=ƌ��gJ�Դ�^�C���p5B[��"q��c^u�ɩ��T���41�'b�;�PMQ��~�z����~VP������m��0D*V+f�!���4{b/�a.���aZ�FS�b�q�.����z�*N�ݓ����5����U]�Ô% T;�i:ͱ%6��s~!�|� �U(���T ��A������omr�pKvqZ�u
�&l⯸Yv/���⑊2�{�C��+�M׻2!�����L0$�)\Tl+'BN��u��С^��c�KP�%������c�\=�즐��9�ܧ��������"��#W��rS��5�i�}�/���܏"��q����3���sJ�ģ@0�|��_y73���7@�b�8?�)��(	��fs�;.�m�h�H�O��aH�c�rHr����ܧ9VB�	�a����n�2�X�DN�W��r�0���ʲγ]���ppN��>G	)� 7D�O�
�X�\�D�|(��ÛT�����	ve�(��a���U9�ĲΩݙNU7 zQō7�\%�-���3��\�,���Jj����rM���5�O�m�p���/9��_o� .���U=H
?`���f��is���"g�\�$��cx�RJ!����������5���Z�@윱��S9]V��܀���9�gw���K���>K� O�{�ء�g㈙S���,I�S��X�y��G�k?��9�r蛆W�8\`�mj�����S�H��\��X� ?pQ����1�����
dO�
%���ۣ�(_���A,6pu+{�Z�تǌ�"\^p-��?`�L�X%d���*\�[\&����43�����m	���H]��:�d2!�/��zd%�8�z,�ʣAwݝJ�Y���vɺZ�2��,��g/��b�ӡ-���eG�<*��J�.(�B�Zl� �i��j&2��)��� ��緽��Qv=��iK��i�ԌE-y����\u�·��q��TI,�"��qۣ�h���$15���Ǎ�f�ҳ�J%B��fK�@�	��n�xA�M^kL�M��즇���]�k�p��~vl!�]$��0�ߞ��cU�v���m�����;�yc0{���1Ed��aTV���'��!���1��+�I?@2�6�\��g.�^�|a��%C7"A6��82�uV�"�J�p9�t�y��W{e��X��UE ��`�0��&G�ky�a��~�ϴ.X��"ٶҎU�KԻMy?�|}� ���#[�m:����A����c��Jlj�}p�9�R�7�nﮧ��ttT!���Z�Rڪ����#7���*�L�W�t:��)@~c������������}!�S�|�	Z��}7�����H0�~���A��Q�`��
�>y������v�<��k�Ge�z������ 0�P��t�"�W�e�|���F�h�ՈA0�o��[J�f��:<��.�>?�_����T���n�Э<��zAg1�EKʢ�l>�ғg�.�}�O|:�K��^TK6|���=q����Dc�4ʅ�Ӽ��/��&��ÄOyܴ�6m���W�������/4����w����K�ry�+Ne`ik�Y�\,�t��	7`�X��(�	�7�NT�3�P��f#Onv4��eJ��&}�=�a�p�;f��_��8)�h��SOL'�9� ��DF>�FA44mu��-��-��1
�k�i/[3�^\VVO��;~YD�g
�%Y�U=~�d�H��x�7wԈ��z?�k�[�� �y7�>F���lqj�V�i�첤/S�RGz�H�;&#|ش��GPƢu���jdZ;A+;`���\��g��A'��(���������V@��i���Ѧ~T�G�0L��-��?@��c���(��V�ٳQ�g�;�D:�j}#�j��j���8�/��h�v�Z�d�ғ���o�q=��[�k�����S.V�Lړ;���:��c��Nj��n�A�"�W��P,���F�����W�vJno�
����X)/`)���~ݪT��A���v������u�3dY(Yµ`���3n�6��͢���y���Sk�
��oT�J��Q��*����D��ZD�},[簄�Fkؖ看���1F��y���)o@#����)%�k��0��9���7���ÜԚ�#�'M��ST�p*�0��h��v�X�~�-�`(��� �'�A�4%w0��s����Y�W��3�L+B@E���@A��{�u-D�3֙:T[���@�iF�%M�����R'�����9�sL��g�>�f#�&��H�R=[�F���)�B�?�-|qFlyu���0����Q�-&P/B�K�K�a�����5䫃���P{�סs�&붠��s�Ϸ���Q��K���Z�5aVg�L-_��j�g�5�9����]p�u��0�}myT�A�l��ټ�"~pH|]���c���o�G p�9�E1�NO0Q�?�]����k�Jڶ���-����x�\�Hؒ�v�Hj:)�C��v�����W ���lߙ�Z;�y�K8�9�����FO���,��r_Ko��sH�4��1��X@��lj<�ݻ�y�"�)�`NPv�T�!V���i�������NÜ��A���Qߑ(�P2�=�#�D�eg� {[���ТqG�B�Uw���I�
�����P7�e�vr;���E����Bb;�#b�W²��V�;Po�?��І5��6yx���=T�!,�b#���f�ΙVܽ���hϫ�����ćj��Cՙ�YO�|��/�,ՙ��eh^)wq��'��d{e1�
�*2W����-�nأ��2I�`��T���݋\��9��� ���c���T�#��,��E�Ϝږ��3�!���{	-mrW��^Z��௢�tz��N�%��!�x`���9��G��5s9�
��8�Tx�E<&�Ԁ��2�H+s8H����}���
�b ��eL�ȵD���B"er Fa)t��u��@aL$'wŋZ=�зA��A�͚)$�1��4�B:i�%��s�VW��Z�elH:Kv�>���6!L�\bq��As|_F�*7��W����H(��u��d�����#�UW~	�\���xU4�Ad��=�]�p8s���D��%�䆐:���� �3�YnF�`; ���^h<Sѳ�9�-*ch�Y�W�����[�x�'G�����{�|(�	~ΰ�.oBf&�,h��� ���[��:t �/�����(8>�Uf�-�� �6+@�V�E`G/瓶̙8�Xq/���9�����x��(���Ʉ) x�j��d�v;��<�G��4
�`�
kb,0Z���·6VK65����S��ohv��3�5�V�vXG�t�v�pyD�^iݖ�i{Q�	l�WqŌ�\B�J_s�>2�?�0�tT�����p�!k�@�S�Wu��e�S�p;P�D��4{���(�[��\Ү��*�B�\z�Q���b~/FP�|+��	/m�*N�'��Q!�R3���d6����o�D�=�������Ey�z��,~aj�4�����3��l:J���)=?�E�EU��a��sG����M���������\��z�s�GW!���_�(��^�P~���26֏�K����T~�kE��,pS��֔���I�DA�i]/L,%^,թUÄiTL�a�h�w���!hD�-�(�J���{��aS��k󃏮Hp$��h�����6�s�M��E��_r� ]�f*���_zc|�^�XlxVHYEB    fa00     8e0�G�3E)n�*�	+���N�᯿h�樉�9s���Pn8Xz'@��^�-�%XKbT����5���&*Y���'�츖 !��SDjޒ4>۟�CӄH�jm���4�Z��b6�H��9���Ô磈W�z���I��c��I�o�/k�Bm�8�\���3<)4�k�:Q���Q�`v�����6�����o�Sq^9+��aD�b�G���͞�M��e�v�hA��0iIP�Z��]k�/)d�ܮ}J�F�4	B��ӱ���~6��E��6G}� Kx<u6 �~�7q���93��@�hg�;M*\�%�D� ���?��X'@�]	�z\FY����ͽB�����ݐ����gO�5�y�X%_���B&�'ʿq��\�OOf�.:��Ù:\O}u�h���@����2K�]A;��Mn�X�� ��Pb�4g�ŌYFb�Nj�+c�=��U��w�DO;���3�7D������ݰ�`͸ē@���crE?*���@S6�U���8D[L}8]ks�fb��o���{4�h�[h��p�9ް+��B��S���O?���b����N��wN��Ɋb_��4N�γ���F���Ii��#Ԅd
��"��*����%��1��p*����Ƴ����پ����͑,eݟ�hO��8߀��צȚ�N�j��U�����m<_����)���иq��Է�;t�vQ�yC.sA�@H]:���d�z�c[�O���ТF{����H����y��;�t��"��/(�9���!5�w��h����_l���6�k=Q�lt��v�&�ٰE��$��}:�Eܮ��cH.L����2^)*Hжd��K�?*���/��v�l��ҲC8�{�H���� �qP19�*�_�!�@�a2�~	RY��"�涣Кԉ��37�� -"9R��^ ���,�t�5��?��lT�9%�r�m<b��T���W��YI8� ���u��AHn.�:VR�nnԀ�īK���<]U�9 �Ui�]éc}��u��_�����٭\d�B[�u�W�����k�����14/K���/EC�����SE����)��]M�I
A@�>�|U�48��!x�2k�$�J��xwY�;fQ���(����f�
���3�_瑑 |�m����k �ק_�w������۰�9�?N�фǈ��t��q[Hf���l��J�U��-eF9�I.��������6�DIH�E�ktq1ޏ��8�mq1�^��{��_;ؐv�Eg�B�)&`\0�\{O"V?�V�R�g�A�ȍ�b @�cQJd�X2Ά��>fjE/��a09��Y�@��Q������^ ���2����k���I��Ъ�4��ը��h��`�9Ls'�D����g�z��z"F���`ļ6h��M�» V%KD�tЫ֕{��N���N@w�+"(D�<j���s�(.Q<x��Ev�V"ʍX �;ec�6�L���#ڈ�'�y�ĊXT�!�~1E:qd�o��}(�C89�,��3��@��.:Z�W��h����S�Ѐ4�i��´g	(��={�d���ACs�pe@��M_�(�S�ؑ��V2�ܜ���J���7�_VB��κ��O�x�����bz�εE�}pb4�2q�~����G�H�Zo�]���S������]�VS��N��֨7^0O�W��n��gz���,'(.����JHyyC�T�Ę��W��Y,}�(�}�{�:� }�i�@�������X���./���ME��8�Ou��&%�3{��z�.�r�袩6Y\o�=,Eƥ�V穿ћ�A����Fփ_�F�aZ��3EƆ�wR5%݆m@=���'�?Y^�fL�a�sp3�b�����B����Ѩ��=��u�^����n7I��Tz��.�xy�l��[�g�32�7�\.�W�)E�Z܎��`�zB�u�py��;�c4�\�w��Q:�s}�)"�Ϯ��F�l�� ����)s�!�w�v��9E���2엠K�w��M�+9N9�%
Z�����#�oA�����vʀ���]�ڙ&:�~�/O��F�f�Ƕ�%�-��U`�H'�j���S-� 朥V�='~�:����y���#䡟�̾����$��#��򳼅<�qO��^PH�"A�IC�I���KU��M�H["g�]�����Q<��=x�Q&����J�oj���m�kcb�R��W�b:�T��Ȟ&��?|�l\�:S&-]��?`�t�.��MXlxVHYEB    fa00    1110w/¨Ci}�ƑpZ�B��z�K�cc�#��y	i��,�dx��G~G�*a}*W��q�sG��E]pj��bԾ��$���s�!���̓�����������w�OF���;�� 
���0rD=�]L�p2M�'��7o�Ā4j��^���[�g�����f/�� P�$>�s[e�<�:�$�� 
�K/5�J�l��/J�?��W��<��0M'���;���_��H+����	t(���m�+9�4f
>=�	'��������S�)�Γ9ark�ժ�p�Ek�$����^AuvSY���t�Y��g�vC����$�3��n'��A�wX�)V!,��Q3�����o����
�*���=iw���[f�d�J�o=��b���(��]����U���bB|��\�;��u�)�<��o"��ψj*������N��"@L9F�21���+@��Hn�m	�G�j����Otm�;��ivaP��Jz���=_`QH�m	�޼��a�V�uw|��M Y���j��T��h7��=��}B��-���M��U5�~c��p1��4���H�����h�w��-[�N5lC^��x�|B:��~渜�˘]9�*��.��g��A�H��Z�$j��Bk9%����ޚ���E��i��!R�A��.���d�vg���[��Sl�>�����W��P�M����į�5��X��(
�iOB.�1^^����M����8��h��֓%�?T��<Z��X��{UF4���]���-�Q�L1$-V ��!�����ifM�0��0����w�,j���4�L�^4�Ga��:�lnK���An[�!8Ԃ��	�_ذ.���!~M,��E;�8�{D��]���{K��w����(�Q��F��Q��Z#s������>���e]%b��K�kz�2k��er�`uT4E���=%Le�5��1��^�������ڠ~e�l���W������u!"8�3�^C�ftt����Hӑ�Ӷ�J2���#���Dq-�c����X������4�]9�b��1���Cv؟Wr�Ԙ�,��%ɹ��Z�"C�S�����w�`S�˜R�$�ޭ��(}�����1�&w��F��?�ko_A�$���f�(~�C��č���Y`�R,�o%�y,��40���oP��.�EC��aE(�!��ಂ,k΅j��`%�����9�����Ĥk���-�����M��oWG$����ύ���g�k�2Ħ�|���g��^��?�-����E�QIZ�(�
!K=?��݃c�T^#�d��%�Ӄ��Z��J2ָ���I$!��BQ����$��K�ĩ�R��=��Tǈ�nX�u�R��� �->��ZYt �uq�@��m�6,�����К��29kx���gN*&v*�q�� �h��k���@�T�]��
芲��������*G��b&H�R��֖���)\_���)-W�����w�
ԉ~1ޑ�&�{B�e�ɡ�.hlH0_��Ҏ��F��M���T�(X`�74�B�&��zC�h��$������M��Fz_Uʉ������@�!k�Y��L���ܝa�"�*T!|f���	��tzO��H��WOC���9�k�K��q��-l�m�_"Jd*nG��}��/X��/�'jH��U�1t|���Q`6;�d �CVpK�3~f���TR�f�읭�d���/iP;�Z���]V!�@�~�X�5Y�T�K�y�~T�Ǚ=��������T�zc��Jo�\�w�c�Uk����Oޑ��ﯕ�U.�L�N���A���'	v�,k�+����%��b.��F�S19f܁�A�h��g�"���e7dǱ=Xr�v�]} ��L���+u��A��6��{fi�Y�� ?9��U���v>`"�����uy�YW;���>�����:m��Ѵ`��f9)�Xvb�;��@k�_�x������k�%�tn�{z3`*��sɅ��Y�i&9����p�%E�r lף2�yc�kIG:B���g�s����mU�O� �|a�����-�P���XX/��H���N"ۏ賦l��N����썃(���s�ifl�R�:ur�9W�tP��6�f�}���155��9�����"}�R�i�*4���ۿ�D@���.b:�V�9>�W2�H�KA���v6��1&K@KA�I$]G�W�Eh���9��k�����j�{���I_u����	��a��_"�f��ȃ�c��Wp��
�`�W2�Y��b=�2�Se$�2B5`���R%[�EzC�ZK��"��F;x�W%2y5�,Ϡf3�z��FvЅ��c���<u�}��� *q�Wα ��@�����W�q0䍨Az�+������ar��[�%#��V�=o<p���P�0�	�<9�VgA�5e��.�Z�P0>�O��>�C��y�OwDŶH��'��i��es:S��l �~�2�~����r�fH�.�/�ov�\	T��, E��O��$�]8�I�q����FQ�7 ���

�� /q*�u��_���,-��)�W����i4r����Ku���"�I�A��[P�z:� ^L55L�\y�����;]�}~-<�����4.�Y�V� ��0�oF=��_�C��k���pO��w�������+��.�U��0�#��!{-$��O�{�#ߤ���o{\bOD��(�h�'{B�!��	���U�^�?&�QmD"�sT�^*�?ǳA��:���	�߆�i
�mQ�HC�Q�:[*E����7Q�L{S��Y��Σ����%[i	�m,����~N�S�(`�FEw�%���	'��~�Ͷ.o'�\�f�EW�/S�u�kоunڦ�>e���4��(��Q������n4���9�����_���X:�^�3XcS{2n�E~���b�Q$g"Hῄ�����m7weV<�����fux(�J�~,>�����S���L,�iv_Ӎ�D$P�x|���d����%���k֨��SL��l=\��iz���U�0����xz�ߛ9#̒n^�;���%�(��A�i�c6� �ֆ����5�XOrL������\ ���BZ�w/Z"}������5y�L ���i>LӨ*<3*����zfL���5�ǔ�^S�s|�ĝx�2��3��q��]�2z�Ιɑ4�_��FiTpk����`�F"�U�XJrJ� 3%�9�'8�w��NO#�R��"�͜`$ȍ(JW �n޾,d�B��C�~��C�Y��S��ʥ�zO4e>��x����[e���s����F4{v��f��8$���P�#j��v������\�c.�/s,���H|�yj���ۦO˻)�'n��'(#��׻��1gn���eM�k^���6M�6(�J��P��.,�Y��~5S�ly_��݁^�t�W��pӱ9�^)H}�^�|�$7Ŭ˭�~�F�]�,}S�^ �l@�������=b���b����\ӕ��U��gb���65$��[�,��8�9�еd��K��V�W����fy��Y?JU���X]Nj, ����͂#�1'%�C��L7��4��&Y�H�,z�����͋�)�b{�Xbi�1T_������#���š��N��K�L�h$W?������Z���c����+�8�~+e��V(Y���<�Fs#P:8�O1��6OK�e-�쨽 �ӭ�B�vwv�Fх��P���&�������Ȥ��.S2�_�ѷ��k�Pz�Bc�\b�"�w�Qk��_�$Ѝ�q�5��r�@U�m[�K��_ƃ!lَM��9&-��T�(%P��Jm樑�``��F��F�Q����T�Jf���϶���<Z�p��4%?�7�hΖ^um�̔UW�Z&��*;�V�}�L>��N����U~;4������A�i�O睧ؠG/6l�^7�T��5O��8|�d*��x�C&��v�})e��l�S>���3-�s��\T���䶻Fa�3�z�����Ȭ~ן�:]��X`ׅ=&�w�	�~e�*V'������雐���߸�6�5���0�ԧm�H���?�@�J�V(����j�M��޺�/�	�M��A�!(-w&���:Y�S���M���e���/#�G����̞ � AjA��c>���(
�6?J��r4w���r�>4!Ϧc��G$�v�����~��z�ʖD
Vܥ��tVAv�d��'A��M߶4vI>�2�4�����b5gi���=M�j=?��M��*�Ķ�,��ke8n�eDj�6I����XlxVHYEB    fa00     ca0s�`��uJ���dM�{Ч�]A~�z��pa��tl����/C�����9ַ�?:�Q|D�S��w��A���|E���A�nI,|�G����f��p����T7��A���8���OV���"���h� I�H �w�>?�fW4㻕�}��+�� �T�{V%zb��oi�U��L?��8���ҙ��z���L��ݯ��^� !�uAS�ߩ�q�pК@����6�� i����AV4#����N�O�'���Y?U79��ժ3!j�B�x�|��y�5j�w�E�"�w�||$����UH��� x��%�?��ǌ��Z��/��&��־�f=�	C�Р����^�H�r�V��T�%�c�M��X��0�3O������w���L�V&"QG���(�KeRE�a��O��Q���	ó������Ȣ���.Vgqi�P�I�כ��a O\}�(�� �9N��T�w<D��Fj���� ��&�s�
o�P1�5�3��!#���Pam�RD�q�q���K�_��^!>)?Q��l��%U���}�:G/���,D!�?��ԃ�H����Gb/��S�
�E0��J�BhU�p�r�NK��8:��

��P�qR�?�:��b����Hikއ����	�)-��/V;�W*ҝ[�Y��D'�@&�u����wuǗ4"�IGX���mן�<�f�9�e�7&��Y?;���U�|��Y�t��\J�u�p-�e���l�v���������G��t�{�{�Kk�%*�M�$�3`G`m�.]}�����(7���G�w	k�T�4lT6� �$W��g9*ؑ�J�g,m��臘|H��H�&y��-� e�r��t��|�4)>����FʂY�[�G`q�j�Ǽ��>��@�U���@>IYht����#�'e�h^��h�P���I#�O���B�J;`C�Lr��W`m�뵇���_��G�d��#���T���Yu_��e���;:�����
4��|��hLL:�7��쐜1h�<�R�h���E��z�R���EU��d��;��?�:��̈��5��V	� ���2)�����Hçi��׌R����0�ώ�b-Ǌ\����3-W��!��L){&� ;�VŋD�ݢ��	C'0�nm�60u#�W!� e��o�Q�O�#a �y�΀7���g�A���#�.�}J�8Iz��g�����(����o��9AhMKH*�ܰ�����#�8�?�?/���(�G��M����hU����L���/o�H�2��*��pC��U���= Aw��ϒ�{�#;�!���pZ*�n�<�L�����X�������ck�!���;��q�1>(�e�w�<"h�����.~��{�?��~�Vgd��ϋ�Յ1S����]�2���J�t�8 ��<����}�u�rW|�$R�4^�)پ���e�B�K��ިx�Ҹ{�ղ���h��i�!�'ls:%���R=�?�Ց�n
��b
IU��,�Z5�<\)dQO��{�ř\�4R��:΅�n�k��o�	S�@i4ē%CQ�~�S�>��8�[��3��;j4JoQ���)/��2p�8�������|�Dv}A�CL�7$�@��W�y�<Z^~����1#��ɇ���7>��[���Z^�w$�0y��_;�҄��9IZ�l��	��~g�s�u�2[�:��$:����ְp_DMih���w�9�^B�rM�i�9W�*�c�����uB%�in	;G�E�|�ɟ�@�~/R�5
�Z���Q�G��/!S4���/��)��r��e@�P���w g�R,�fқ�����ƎZfoX��pD���W�}���b���h�M0��B'U�����K��7�@f��~DU<]8l-��҃�gx1D��} :P^_�2�48qr|�}�Z��q(��;"gR>'Gu�Ѧ���UJ��m��T��`	9�����o����^ j	d#J�{�����ԝ����S�V7�F�R����^��Ӄuq�A�3�����W�[����.���|8�C�j�e����+�*�X�d��ܳ��^t�<����e�����<1�f}��~6����Շ����[�{[`���@��S"����⸅��AC�e�����W��B�0i�.Њ�96��,�A���c��m���_ζ_��Y� �QFs�.��A,��W���r"��que��»r�����z���$aJ����_��������D��"�j�T�s��Q�Oe5/;r
��S���o��{JI2�_.짫6���x���{��in�(����g��4B�(|���E?H�_���g�8�zHT�6|p����Dd�������ʌ�9/|�M��R�}���x;�5 ���,6��P��s_Y��� �-8
����͐�aV���R�WI'��JdmtWo��=�I�9Џ���%������n��������%�rpR��-V��!�i��,���Ĉf��5�v�G�(�G��G�
KA{� �x���g��,�{��*�`ǿ��j����z�{Dj37��[�@��)Y����
N�4�8>�f��e̠��s���d�����0b��<M�vz�$Ss��g��~���"���ψ�+aN�$�s�������΍�q�(�0��W�����KN��8�@wo�q�ql�����C�F��!2ҭ�̇dʇ��X���῀����mzzW��'�"��-U-�*D�g���N�����o�Ĺ�d��C繽'kq�M� BgT_��-����=��K��=}�0�b݈%SQ5���kBk�����T�Oӥ�������$��n�BNC�=��k�1[gv��in��r<�즾R�ה#�#wϙ�����{kUb��M��u1:��P�uh����G���g�y�*���`i�y��+����f���)2�Dc�n�Yt[���&�SѲ�`T�{�xW�4�THйT2 5׬��:�w�|���+Y�����'����K2�=���GzV@a�1 ��[jA]��aj�^]_��Ã	6_e��Nj�����M��}��7A�QMr�q � AuYπoΣ�9���N3$��֘�7�|�\��qCf�Ln�4�k8w�HC\�;����fhD�tԒ	��B��Zu�<��9���.��$V�����~��4��G��2�mS�2v?D�����XlxVHYEB    fa00     3f0y_m�	�RsW �h��p��F��˓X@��������Q��
Zx)���1�{�rݝvݳ����I�}�1�� qy,��G�;B�=@~?������8֠�6J1��sY{� �E}��w_
o�G�dp ����zH=�=>YF��!�k8c/�Z�w�Ngf�D�G��́d��U�m�yͻ��U�˒i����ض= |�h�Ϋj���f��x�I���4^��H�)6[,��BU;-N^Y�b��c�����^IN�P^�G��J\�v^Ѡ�]Y����/���&���S��ߌP�RFc��>|`��A�˿�1�xġ?�������0�@���
�-�	�DM{�#�Z&/؍&��p��y��!��t'LxS�Q�&C�m�N"�ހ~׉c��fڨ��d7�ڍ@��֚_�^�EI�z�q����nZ��-��k2cw��c �(�`� *L���aZ����U���Q ���tu����\P.l�
����Y�z<4uq!5CTu���{/r��l-{1.16�Q7qfw�����0G���N���3�c�^lD�~H*�b�������5�9��g{_:��Wٛ���MĪ�UIH����9'N��	K[ϐ�sX�j	I'H.6�=C'��.pD]��$��!+�2�֨m�쳚��!�ik�܆��f�<�D���R�{g=(	�Dp�d6,|2�7���t`��g�ձ%�8$˫�g�g�8���.�Ԣ3]�BV��ZO��=q�q��MIܻ�畴U�͕�̖�ԒMq p*_�0�ws��-;kŊS����Ǵ!�6ɩ�&�`�5l-��8r_'}�[�Nx�d��@�)$�1
"<��s��x��sx	�ĻxV"αǓz~�(��ql4����9�?���k���1X}����j�̤~ΙSz�	�	�aAn#嫈KO��Hߜ�g��,�?�#�8�P�u�9�|����!�L1Gl�D�O�]�;k�0�z,��$^�m�a�U�vwX!R^gt}�$�-XlxVHYEB    8096     b20e�c0�tcL���#u��_3)97͘�����"��K!���'!���uҗ�zv!�#�V����l�炋����?��8��k�꼦*��o+��(�C�X�đi�<|���4!�J�F�t�x��!Ɍ�'A�rJWV��/��sgǑ]7��I�zY��d5i�&C1Hi:��Y3�qɮ�A��SD��S�� ,��G��E�Y��g�i�)Pɱ<;N��h�5e��;�V��<���Ttk�2�
~y�&� ���An��vc��PG�)ɨ�G^��9m@M�a����CrIk��9�^���]�ЌC�#@�y�L��`\��#�'�ɕYa*�bQ眏 "�����df)�����^���Ik�.a=�#��C8w_6���8�uF�]w,���<<���8�W��!�v���\.�z�<L�ey����h��P휺����;f<��׍:ʷI��sxs���<�d��a:kA0F��r [�#U��b��WVšG^�C���v��� ���R��������+bN���]���۔���?�gV�f�$�yo��f�Y8��]��w)�L���'@ڟÝ��G�D����Ӵl^(B~�ó�>�������嶓���lV���%��|x�}AXW�?��	�G�D����{v`��p���Ґ�hY�[�_�=:)(/��F�5P��gsD��P�ڹaET�����#�}z���Q��#{-�*���6'�|N-O�O�s�'{a���཰zTR���!�Zd*<�>��@S4>C"���g�*��j���V��t\��Ϩ��k�3�:T�A��(�ҨϠ�Ra��0��`��J�"��Ylif)�W�Џ�=
�r�X����ʵ`�zf$����z�Vf{Β����?�R���͛����j��r��{�D���GDcah��a(Xd�Aˣ����8Jj�4�]s���5`O����m�b͔�ΌΙ4dh%��٦�kk��։���Ƙ�������q+h �?��m�p��c߁�%�����րe���`�����ޑmf ���L:.�p�#�Q��94m�W�>��Nj3r��5�i��we�&�G�?���	����Аe�����&�L	��̕�#I<L���H���E_�)Mi/g��������.��
��9dp�v�ѽ?fI.".3�Ye	�ۡɢ��eƺ>�4�D�m��j9��i7����?�4 ����8ٲ[����x纙!R"�,F��*�.�yO�7&��AZH��H��G����IZ[n��2�_�?:3�6����E����Ťj�{U
��V|%f��' o�_�*�~M5c�?�M�D{w)7wu4��v]�斪	%�
] �s����s%Sm� ��D����Z���g�ut,Me~Bq&"���R�4t6ǲ+��Fg�����o~D]�.�WfŦz���K�PzMZ���%��U=}���H��Taԉ:��2�*-c�`$� e�^�?�3��p	�K&.%�:$����)d�k�.�:�ٙ�_V�p	���^�JWg��˧Wha)8P���{k�س BN�C���`+�I|j{X*hH�$�	w~�![�P(q��!��_����ߧ �(}���5?O�bT�ACE�\kЦژ4�:�������I�ؓ��M��Y����ȍ�ϗ��孬�Zx�Ʒ��}��K5�d�'X�)�� �VGy���My?j�����k}��Kk�Y�b24'��S�E�U�k鰬MsAD;�R��Rl��9����D�幌� �_�MD8�z*Ǒ��~&���]o�)��^�`x�U��GnaCS%�0�mI<|��޿KyY�7���&5��7ői�Ƿ1���S�y`ظ����ʳQ�)��e��	���~���)�E��{�7�j���Lى���=���$�UZ�?���j[�VZ�>&��>�W�[��J5�u�tm8ۨx�1�1��_%nC�����u���髠�J]=�kjf�e�Ͷ)�g�G����n���O�Af�|V�9�%&N���{�c���Q�P�R�\d쿲u=�Xr�ϧ&�S�����p(�4tn�Y
�M�����!���m�c�>�rS�.�@������S���3������y/��S@�L�c����xW���` �q�������ؘ��E�s�z��g�6��.'��Ġ���##{�/U���x���l��jG�P��N���<3Hj��(�,Gk���1U'��,lP#������%<NL�`Z}k����}�����~��+גdX�k��c/���N�0���2�A�"H	{�ů ���*��t��B�����p��-ԛWι���$��f��91�tEQ��?�ܶBQg:uar������Q7�߿ss���[�����e����7%U�y�#��v��X���"($Ц�i-3�������'��FV6�:�4�{A?(W��0�e��hz=O��8���&�������]jq��`M�l��K�"p�46G*�����V)�f������7��M!n�P�K�w��h�&�Y�ܗܕ&�n������0�����j�A�8L#�;/�n���go�`� �1i	�[��ǒ��=�~�f_�J�9[�T|�Jn���^��� �I�3m��|�E2����<@���T��DW��%�S�����h���^��9＀}�-�$z{�ִ�"�e 8}O��D����B�p�0�t��PY�x�e���
�2��#o�#�K���ȥ����T;�-m�Fa��zv�۝�%�5 �����