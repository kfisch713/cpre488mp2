XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��DN�lD/�ʛ�� ��z�������܋��w���x6�qv%ne;��d|k�\j�X#�?o����AR�~T�D��;S"�>ǿ�?�V���}�g;���6z�dP�b�"b����x�O�����}��@�]0��[�f��aX+�f��[o
����
"`�~��A�T�v'x
.��.��s�rhK��{c�>	qi�VT��4 hc�}��$�ݫ�}55䫉�%v��+��B����|��/�,(=��WTl>T��ѽ��'�l(�D����"i5q!P��뭘�p��&`A���ڊ��͉�*2�m�_PݵY�z�9�Ძ4�P�.���P��N4T���d�Qd#����0��,WO�iI
J�zǝ\J�pK{�G�����q��d	O"}2�ス�Ұi�R����{��AIW|׍݂U�D��v�L$��n���1u�>WE�'��d��/zŃi"F�R�J:vP���B�V��2���h�����m��;S�B��� /�K|�� $�8�|��u����AV�4`�r۝NJ�Ȯ���̩������#0[؃6��XZ �'�Z�ゼ�m��Q�Nv�i����*_����録A_�YF��!���	�,��YA��.Jg�2�ڞd����K$�A:NY�ehd��c��(����cfӊ�oڳ�fSy��4�������$�!<�́�V+8<�mm��#e���倴�����Z�`d�%��Я4p
�;@���ls�N���<mXlxVHYEB    1a34     990��%6$���'�Z���� ��.'�_C7ڢ�	Z&���':u��V1;A'�V�9����*��=�j�
�\��V����lɨ��_��t���Ȇq`ah�m:�d�o �ظ<�k��d*Hݛ�rMN�ŋ�O � �e�G\b���qU�f�N�;n	�\�
g���͔�*�[�;���1�ڍKn1&Yԟ�Nx�>�\�T�6�m,[�Վ]g�e鳈���,7���(�黾̂���']UV����q�� }+o=E�ȭ��$�7�~�oyQ>ϻ�=��"��8�u�R7x����c�pAtB�z�Z�	��f'�B-����|x:��ƹ�o�i^�@��*��J	kWy����ӡ��I���_�ʖ��Ɠ���O5d�J
b�O��*L�����o���_��E���`A�~�SH�רb��ƈ!m�Z�=\5TK�N����T~��D�HBJ ��o�d�v�y��.k��!�b��!�A:��.���W�n��	$>��b���av8;~)H���K���A	&�{t:�a���:��aS�)5�`�W�	�yT,��c�`����b�¨�`��4���!�x ��]'5�7�l�P�C�����o���p~�����ZD�㔞�@8^M����7���@��O��^�B���1�T�䐣n�s��a�|i�&��������7Y�J�z��q�b+_�|��d} ��"�%I��:X��)�P1lY^���է����8L�Pe�L9x���	NZ�Dfc�a���X)n7�5�8��5�D� מ�7RW>F���q�3��Aޔ�fpc
>�6iAvr�P?�"��5��| R�#���)���-�H`��Ξ�b-q��Kk�h�j_����A��@�8cA��p}ex�y��'�v3�6c(��T���i�q�����N
���f��?��)����eIąI ӛ2T������0Օ�U@>���39��Bǥ�Sq
��k{-|�m��$8(o�����N�ͥ�.Cƪr�Mb�tw/�� �z�X�t�dn|��i>��c��E䢔�n�r�*]��$�K����Τ�c�w#��>y���$Ir8��?���Ɖ��7��6G=�JxF7�؀P����]�HxL�{�9���j��$
��3>�nt%�K�)�]�G�R#O�c�QV�dHN4Q?E:��3�H��;�l<
�0�$�^��|��L!*�C��fŎq�5�XQ� �?�v��Fr�x����3���̷�6�(��W�%�裈+�ª1��Y�&���r�w�v�7����]��ڡL�������m�]�J�T?(���1�U��C��-?'6G�ʈ���z	�N�v���Q�������l�v��ڄhzǯ�_���A5�ô`�Ld�:�v�IR(NCw��J�#,�2���a�<a�5�:=�q�W XZo��ȹ�N��A���\��\'r���a�lҸt$L�
���%�)�Bu����Q>�ta��Ԛ�N��i�cT��(jCu� �Ƽ��ݺ��s�K@V����wS���XI5��^􃄰!�6K[Fgǵ^� �Ƿ�1���Gft=���NHI/<μL]��}VE�\�`7�[�UOZ��~��$ࠆ^�S��cv�A�����S8	�r�Ҿ�Y�ޠj��;
_��3bg���'���ѡ0�Y�������h?��S����K�	��Q}S"� yjC��s������=c8g��@d��ת�,wy�Fy:���Cf4��.7���(o�5��QOmHc]��3'�8b�RG6��:�>�q��]����ɡ$n�Ȱ��z�3�ji	������/�mA3��Ab�~����KX*�WE�;��gݴ�X�����Ax�����e�:,�E]W���K�=�@���f�j|�ƄT���U��|��:��w��	�J�s~ou�P@�n&�����Ԇ�t��-15r��������%ZwI���D��'��M�A��:�.�V�U�l��yo��oKr=g�s~�e Ԭ� ,sfL7�ku��#^4UKֈ	����U��cö��z2�Yb�Mc�|0��� 3H�|�R�h�C��9ݍ�Ay��A�Ñ�8��	�imv��s��Z��veEF�Û6�u���vQ�$}LeAA��4	=>�!�}�D�f���� d,L�cY���p�d��U�T�:&X�����}͕����5�si��K"�}�ĺ9�6�N��.����d�j{Ff@��i�H*9�ӭ���K�S�1E��U[�65~Z�m式-�
��a�~M{h�ES�f����~S�Ϟs/OȞ�\�T&���Ǡ��n|`��[�RU��A����J��?IF�f�6gX�
�	D�צ���c����|V�E�6ńh:�^����K�