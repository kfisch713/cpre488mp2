XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����As�X��5q �?��{�!�za�A�t#/�ZR
z�)�L1�vf��xmy��9������(a}dnȆ t:�r��+>ܡ�q�8��\�}��%Er��vY�hۈ�y-�);L. {ɠOx��}�����t�VZB������R�Gq����#̹�K
�4��j T��!�$���̢��B7�"t�)X�H�G#��v���������r�8��ɞࣻ�Nmi��������������0˘2ı��Y�m�<L)�C���3v}g��=KZ�򇞛���8�\
3.��qS\(�
�YK��"B̔���4h�F9ӧ��C���%k���tU�k��{&t�,���!�� "�.	��{�b>���C\�=؀���>�-闵T��x��>��ɭ[����,�AO��/�q�UC�y-ԏ!-6Zx��`c��{��{�@�I?���BR��6�<튜7�ngK�*�q�dP�� ��Fj�*mYi
K�3�ɅV��;J��f�Y�M��5����|A2y��\��,N�>�d9> "��Eş(�u����v-IOV��w�9sH�8�!��-/[�>S�������3����+�=.�cp���ճˊM<7�Ъ�p��ido�ϟ�w5cc8N�ԛ�z*y7�w�(�1w꧹�����9��U= e$2�W�,Q[��6� �]h�	W	�E���g*�V�=��ƀG8n�.�Pz��{�ݏ�>���l�yPjxL�~jᱜ�F1J_�q?�4��ćXlxVHYEB     e07     680����\Ơ���n��|�Km�8��� �Z��A��ޱj]������Av|�|b0W'�'�v����6�S�#�I ���Ek�ā��Hb�ΥOS�$����z���X@��̾T�:�KwV$&[�oksifC��<��+m��ƧH2ɤrk���k�TD�)�oia��-+�}J��<��C��3�����:�?@R&(I�[0�>�V]�Xtz�`闤\r#&+���3�&�H��r����=h.˳�_eG]2�R��*ȅ;Gbm6�
����OK�T(�=�Y���N�L�Q�z:�MB����\nErʰ�&J�`į���A�;��f��W�f�,���I8�ޚ@��J�	������	b�*�y@cg�˃-�F!{H8���+��$���i���d(�������ׯWh2�ySk#��y�K]�#q@9�؀B;1#���t-�zv�6=�>��|�xO7���J�#�++��olO�%�gt1'3i�Z���:�Ҋ��-
���⟼��S��Y� �K�g�f�9���Qt�
\+���^�ߏA#1��˖��}K�H��.��,�`���G�6ieAC�@�'����%��z
F�@�AIV� ?�������N�8D�d)�)ZnZ�]�Li4nJ�(<qL�e1�jŘ����,.����KG����9ĺ?=g���:_)���Lz,�~SG[eY�=�F*���>�R
���yV�[�1���F����x���l���Z�/��h/�j�vD(��=8T$����L�GC�d0H�
t�aǼQ���푵N�`��'���,!�# �f�0�P�BڕԤ��ړ�j��i�m�.b�UT��s��ڑ�x�|��^���� �鯮�P����b����8Wxg��m�R�i������=\�D�ƈ$��l���`�'ɠ�-��'��jT'-3�� �{�:��6C�(�tL��-�����G�258�B�s�THB�-,;�H��	�Z������؀�ڐ܊���M�r=R�����)'����F*瀶a�����T��g!^�~�ڌ�f���DP9%�M�K�fq8v��3
	��\���hou�f��o�>vw�\`�8�Z������K���*�[oVÈd9�?�Y�i�`��B���w�Ex�kNdNZ�ؚ?*.c�R��H�p�m��&��ZC������S���z8�c,��Q�4�Q�n�C���&]da{&��:o%fZY~��٠��D�v�a���I6��W�Ziy�����N�L��w5�?��j0���,JM�8Ax�m�7���ϔ
�0��/u�@�ĞJ������u��1_��'Vn���K�s*��gն�h�퉸d�'0�)�25�<=m����͙����:WzpE$�C�QH����)"b+C@�湠����K?F)%1�]���@��	M�Ew��,׎o�2�}�P�<�W��UR�۸�k7 �#yAZA+l��*� 2���Yb�;�x�%g��`8GQ:�� �G�#���BU��\����ԝ`��,�1a��P�� �Y�+��g�=����p��qH#�F]�ɭ΃�Dt���O�niT5n����1��w˾ދ7~_��ED-�e�d��O���Qb;eS����1	�kr}�a_$g}ӏڐZ�