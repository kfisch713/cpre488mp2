XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5X��ـ��дf��Z�2G�Q�K�CbeO�f� R��V�Wt?D��Y�R�w�Po��D��VPA\�X	�j� �%�1��G.�P�A��$�]������@A0ޅ�K߉�~�����ϊrK�\�̻9��Q�����?0�v�� �=�aw��L�x��t,����ic�m���4��~��?�-����<#ȁ[��G�YH�U-���)}��~�ꤨb��ɧ�@�8�o�'h��2p���XB-�L�T�t+���!��Fi��4�"�d��@��u�����c��	�p�C̍�S;�u��C���Y��`�a+�lO)?�x��1�1a�scw�}�T�-)yDkW��q�;����v� �����ӑ��<��_�;��O[�%̀g��X;R,�J�*~����C|w��l9/����-��)v�KM��)u�K�i��|�^� !%VeX�l���=ع`^��#���ST+irr�0U,�y���/6�wU|�1\�x��=�T$2��~
>�#�ӔŜ�v��.,%G�qe��2{ \B�[����1p1���m�<����s���0�P��9Ҏ+R?ٓ��#t�GZw.s���a}�:������y<-�#��u��u��*�/�'����)+��$�5R�6]�ղ�� �ǄM�[7 Lȴ�э-S�AH0�:��B8�Z�v��y�߸y<�#F�0���������#���2f-(�*`O�������������8ϱ��XlxVHYEB    925c    1a60>M'N�+����a$l�m��7]x<՛{f%C�g�.Z����r����3D���&�W} �%߭Y[�����9/͜k;�NR��-c��>�z��~s�G$;���6�tr���kq�� ���{��0몚���s��)���D�[�ͽ��R/���TO-�t��Je�~��ǓΌ	��%%;ʝR�.�U�8��$���S��P�7Ӄ���!���CHN�g�ډS�M�C�_��->65˨������]��F���I��
T�gʜ������r�^�X�gF끻� ���:�Q��!��S7�
�H&A�Q?>�<�7��`��o-��̇'�"�o�B���!U����%N�8���ݲ`W��4G=L�ӽĉ�%��UxШ�8����P6F��K�1P�@�|��:�u���V�j�<Rw���
P�%�k��o(5vӵ+���I��;���X�M�@P�|3Jq⏶� x9"�c�#�H� N2xx�?YLM8j�K�ڽ*�DQ�D�=��Ĭ�5J�rƯ���3�5 �w��C��&�Qz!sd=�����3���<8�)�N�1KI���n�@�H�G(C�nU}�uE����\��q�L�3��43���ZQ:R,�H):A=bדs�(29N�۞�)�m�j��~G�.j�j�SCO!XU&n�0َԩO��lYt	ڄ���՗7�(vR��a� �Bd�������vX#b|�s,h�L �Tw��L��飶���A8���j27�&REÒd�ρ.��TK��Ww�V����j��O�2ہ)D�o�� 
��1����w,�� �h�N��}X��.'z�c9���s�[�Yxp\�`c`��K\^�֘��NY�_��z��������W�9�M�����6��c�BMHEE�n��>��I�~�o�����`�N��k@�͗[>�:�ߜϷ���E�Z\��n�ϑ1��',���k����lܯ|�.l)s`�+^Nh�F�&e�J]��ȡ�c��Z)�����@t�Vƶ�c|�t�T<�Gfy	�F\ש�2EцYV&}��s��.uj���?���v���j�v5�1A�_M-"!�0Ha�-r�u!=)Z�gFWR��$MPy�Q�=^3\ x!�w���b�.:�0�SE�E�M(�2�X�?���E�f#P�"� Z�?<���9O�b�J&x����8KG킐Q������׃���m/�47�3����:������*����'�;ր��-S	����U|P1�mz�-�N�γ��D�L� ]N�o��y!��j��2To�"�N�#gG-DL�R�I�����Z9ݭK@����4�C_���I,�q�)���#0�(�@b ��#�&0�&�z)�|�	i�5�^��=N&����/������hͨj5x���J�neF��J�+e����v�<�SJ>'��V�fJ'�] B��y5P�i���A`�c^�[���v������h�@�M���/ ��� f�t�Â��\���>�Ve ~H�/�:����k�<��a'N%�񊳅p�CIO�l�ԏ9�V��ן��2��tC�,�;MΦJ��]� ��ce�>P��" �8&5�'��O𕼳��g��"���Q@�?���]����`،�������],�gK�P {?�]�˅�%j��Tl��6�����䟞�Le����s#��HMm���L�u䓜��n�b�q�Li��;�֒�v���ew��DhGL� ��{}f����-���}�pY঻�̑��SB��Q�[�!�	(�6�o��m&�hd��G�H�T��������9S�%0�Z���*���X��NR&��S�6�q�:A����.�ϝ� ���J��&,�	Z��>ٞ)�Ŝ힢2�D 9Hwo4�G&�5�>-2v5�"���P��Ж�����'�w�q��К,Ј��S.bQ�� �\daT�3�Z�ʞkq
��~J���ք|⚃�+AU��x�#�`6l�E�z~e��Fze��<s��L}�ә���"�p"yw��� Ti5������w "�Q� ��'���5�B�����`6'���p��7c�9�:��i�T\JxQP��hr�M���.�]�g��L�)$�+�MɸD�z?�=҅:+\`����'�>%�s�bO��.���M�vH��3�C8����������+���EGP��@n
$���V4��*�,Ch�\[PjB S5Z��W�-����fD` �n>7�_�{��&�b�k�cJ��lC�+g�Zvf�U��j�i�B~��$j/�mS�p�<��PT�d��|��~��/mi1��M������bW���Ɣo�j�q!n�����kHO�L�zPs?cyFbI�w� v�����U��t �g:G����9�}�T�7�PR t�����]�v��1"�:�/փ��i����J��DXtl~��}���+/�|�}9����EU^�ꯢ�Z�ϲ��+Unu#[:À�ɭ��7�o��C���H��y��r��C�0#�P<�Fh�����m#oag��e��$D״3|��l��E�WQQ�۱t��<���^��
;m��f�Q�U?��|�E��(@�����ZJ~��vU�����g���H+nT[�zD4�N��o��;�zII��zxbH�.����z�	~�+���p6V
�4be�4����E?�bSc�b��pNE�@Զmd�-�������]�?�Pb&����m �H�w��6U*q�h�Rp#�pr�.�_ #���y��@�1��`�x7:Fv�+��6�;!ة쥄���|���C��֎�ϔ� �:��ɀ�
�k�(}�<�3D��mi�ǧҹ ž��w1�^-3�]A�dP#��<{@KI�=���z�F�;��F�+���~�*Z��oBve�`h�'Z�)ه���I=�v�)�wgm1<Qp�Í��i����(H�w���݈�&��ȡÉ��E4����/� ��~'f�'V)h'kv_Tu���̴�a�������g 3��!\�S5�x�JN���n��5����R%���P����k�ۯ�)�^?�G�ht�o����p��Q�̩s��z�S���$)/G�sH5�?�L�wo|��6:��J�w�F����{t�7sIe�QN.��T���Yv���z\ �5���u	��(�5i>�8lX�U�6X��6��A�v�t�jM5�A.kU��RC���+>o� ��C@�p��Cb��fpއ�l���F-���b+w��d��P�n�˵[�����[wf^�\�Yڲ�2�Y"d��k?�M��:��� �m|���5f��Ě�gۊ�v��RPKe��u�oN���CܷL�v�mA���ɮ3�}���j�|�4@9�-���Kq�k�e֫d��el�#�����������@���Ѻ:��}Z�>�["���_֝��(}�U�T��s�]$����������O�WN��h���@x3��S"s���=��Ei,��2*�!Kh��Mm�HN�m��=��_��:��T��
����o�J��W��όR�ui�t�X��yM�-j��OI�V	=���I��dc���`�e�iU��KO�_��<Β>��ƷR7�&@�8�.�&%�i-���?�9a�@H�-����ҋD9�F���ÍGg&8̵�D���,b*^AZ�4V�`�*|�?��P�ׇGW��><GThj�ʌ����	
��\2Y�{�nr��<�h�&˶�rk�M*�:.��&h {�%��1[����w�o�͏�3ͤ�߁�K���8\��Ǉ����M?
�C�������h�ٮ,nOØ�D��#�rt?�$Z��	�#�wK�Ec% ��O�8ؚK}�8gz���f
ɳ$xR3c�
%C�2���j.������V��:���*��r�[�B�CО����D|w�W�&�ח��;f�'[f�j�w:��n�Pt+����bb�	W��ZZ���K�d�[��@ယ@�z7��;A��:;��!��amW���N�|l�}U���;���a������`�I�	�����	^J;��E4��v���e�1bI-���A�4�ǝ1 �؄H�Y�}�\Rj�`86�O��ƶ���ȭ-+��<�b��>(sO�� ������E^�ʯ������7�m4���#���Jo��9D9��H�`)9�7�I
��%�t��/`Z�t��+�H���z�̟DYh�f�/(n[��A�p�|�
@�g|}�IW����Y�_G�ӓ�}�Ț�,B�]1j[�^=���s%�◅f���ʹ���aP�мcփL���?*E��X������{m|!V�c������&P���&��m4��"���C4nɂ��""�+����V�r�1m �:";�S�8j��Ԙ;��Ƨr��G����X;L��兒������'���)u��m�I����<�F�W|Yg����{��M�  kP�*��1�!L�Ƿ�
�|aE�wR80|�l��؂�r��|�3e{��A"����n�+�Ywa�,�����~�	�Bw��4�y����(�
�9\D�=�Hd�m>���՛3}�>��":�����Ҷ~�eZ����$�:K�/HR��)E3�����n�6wTfx�����{�p}=	�&g|�x6�.H�z�(�kŧ�l�h: ��(ڪC�Q�l5�z+��hFǥ��#R�&wf%B�2��{�wJ�B��1ak�&��f���QK���9�D����hk�X^�S�n��md�;R5Ȭ��F�W��@��M���Yz�B^�i��(�4ˬ�V{�ꑾSw3#X�W<���������u�6�_*�j�p#�K�	~9ʖ��E��|; _#,(�iY�=�j�@s�8P
�T~jjP{�����ѝ�]R3>|	�wg�&t�X����CD�}U}x�:����@%��J���a��9�� ��������,j���VÉ�&`[Po��(���쎝.����̦���\Qg�y���NE�̵Ď\;�"l�!��]PȀ�Di13�X~�Mk�4�.��^���{Vz��ѷw����Q�%h��kL�"_P	���c>)���
k�EI��qQ��Gݏ�.��#��F�;&go��fQ��5�zЬ'r`bO�e�z�H�b0�g �J�cHL������
{��]�%��!3���� �lC���ו��w��]��y�/>��V��w[��{CL���`mXĪ��e�T��_*�jk�H��{�#P�5ܫ�v鉶�M
�K�p�2�K��#N��.].iw<������?V��u)̫?�-(<�Am�QޮD��O����S�����%�9�O�����*� �a�r�����:se�ɲ�icG�?c;��������l���$��k�bˡy8��\��`�xS(�A�����N`�ގ�G��)l�,&ãY�j���Mr�_\疶e���+�}���F��F(j14'Av@h2���=}p|�݂y�`�W��V���K���s��Z�V�N�"�f �d6�"<�T�c�ս-wYm���Dգ����TaH��Q�Ӽ���6�4��f~��`�>��p��8�(vA%S�.�I�ڹ���qJ���ɢI���}AgG���{��9�C۟�[s����������ŻwVK�w{�(�����E�O�x�!�g,I�'�f����U��ǆ_dQ6oD��3��կ?��SWr�i���gz�H	}���E�|s�|*�F��Xa֝A�ɚ�'�|���æ饗a�B��(��&�(ZHo}��"iJ��`ǳ��^ e`�Q��IE+>�E/���ȹ� ��A��MM������L_���YF/	�0�$�+��%;��Q�H3G0n��a�*�EOٌv�1��͎�?` �ϋ�^�B
�x����쵝���9O�]+��ѣ�oVnU��f��y�b�ޣ�_ӎ>v)܅,C���ή_k�x�um��+���W�)��_S��i�`��?�s���ed]��G^�>�}U�a�@�1cu|Ӫ�06����7��g�V��B#���M}6���,�d�[)��JP����4�giӺ0����W_*>_�ƃC�J*:�0��>-T�n����p!A�7��u�w�BIf8ͪ,��&�P��a�����utͻ2�)�vi
 *n���	O�-�L����_��%w��'�- �V6H�i��XԏTͺ�.��������p��}�#Z���b� XH���"��g~��vQ�t=�ԍ�Z�耢M:�EPK� ��>hb�.�Gq��{x�j�d�\^��o|�w (��ETy���p5��lsR�K��W��n�	�R#d���Bڨd���=�g�T������)7<��!q�-�w�̞ý �f�)T���ol}����v&?Z��L�Q�b�=�_� \J) 
%��0ڴ5t1n�X��C�#�r��NC��IS�{�7t��l�ѻ�������b��ݳ(`�M@�ѫ�1�蠅�7��ƙ��a��蟠ꬢgع�i8���m �ԷV5��0���|��B�,�iЅ�����i� �5;vx�g�~ё��r hxA�� "�(�yh-��i�V����T�&���ݫ�	j�?�