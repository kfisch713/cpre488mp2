XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$�n�2"sЖ*Sv�l�����/��'�E�2�&��ޭ�zE��lb��tN`���N.����;bX*1�z��-�ۍ�����!�J�׾,�W�16%�n�Q���a/�jFHV�v�:i3��}~�Idt^?~�?�柞G�A�!Jw�6?�zұ����K�Q��&O��	��g�*bo�zY��YLF崰 �d}�m�
���B������	$���*O]VI���yG�.SR$r��<g��vu�<�FM ��0O�g���>�\��	�7òp�b��CD��Q?���%�9h�Q(ຜ�0T�	i�ڭ�	-M.��T'4[���GϹn���٧P�kn�_S
Z'^����QE�}|C'���
���K�椓�.�wBQ�k`4٠L�N���MZ��K�4��Kp1!�Ep:g�n�臂c�����'��Q|��ϩ���o S'ՠ�[v�5�}T@1�j��4�T6v� ����8Ԓ����ԯ�p�{��_8L��.3�����<|e.����(�&2D/F[�S?B���_���?��W���k�Z����������E�H�q��e��`}h�c��������/���66wT�K��| }���	�3Ý3�4����aa
�n
�H��;�A 3��p�����[a�m%����eِJ�!wc��{�]�,)����̶�z޳&�f�����ׇ(��P�6ō}!����Rve�"������O�y�Pg�zrz���XlxVHYEB    5d54    14e0>S�:�!Х�H 
�{�a,"��D�ge��,��u�]�f|� C� �<��-��!�.�*���	��gHFa���S(&{�K�א��𚶱�0{6�b�@��hTS,.�Z�^�uK�h �	*�w����r�m�l����'�'�,ň���Av����({��$����ɻ̩���@a�#|����`��^�f]Ę��d��S\�ۗ�#z�3E������0n%��Z؄�w�1EJ3���W�~�4G+bǮ�LOK�P���!��%J�J�Q���M�F�o�g����BW8��[ݩ�O!��k��� a֕�V:~�B�e��uޣ>�����CPh1Vzc��'�/�v[�l�� �&6�o�S��ƌ�9��7z��HM�����$O"� 4e�I�z'v��ᆮ���6.�oE6�lؿ�'�� ����ð.���(��q�5����#�6Z���-%�ۓ�Y�p"�MJ̄���,�E���)ӎ7 �U!�1�i��ux���A��׬��s��O����G��ꤙ���	��w>c��RC����D27�JzW���
�����k�?���� �� ��
�|��V~���z��u7�\0<�)Ҳ;ֈ��i��5[�U�9���j,k� BN��:��±7�,�H 9z��	����w���W�DݾW��%-�n�ɶ�
���	��J�=D�	1�M�ȿ�D�d��{d�b�l�(��VBc����Gb> ��&��O�@|~��G��޼\T����Ub8S����o�`L�ܖ�%o�,xZ9JF�@�k�/��̴G"�(u����"��������h��Iꉳ������p��R �%�zpR��m �u�_1􍪚����ܐH	/�:VAa�{��.��YQϣ�:�n���0���N/��P��ˁ�%�V��(���{�zDD*���|����;N]�s��g4I���S����WɑVX>9D��4Ŕ��tX�*�Q�vҚfcvy��c̩Y��ub��a3T��nJ���<�&�0�����4�l8�\�Z�8��c�7W���~aD�N�:�u;�hj�D�qO9/��E��FA�H��P�Y
V��}�o�i�#R/��e�'��a��n5oՆ(BE����H�c�H���373�TG]�T�Xp_�?��Z�"�Dh�hh���
�֙��:��ஂ�>�!�&�uUm	pC<f�O��1����H�c#9?�X��o���o�_����ܥ<��K�	M�ov"�����:�^�C�\�	:�������[�D9rq�V�;a��s��.������=�s2��b������9��e���;��0Q�[Qp��a�	8Jn$�Q1�Q*�?�ݯ�PWL%���\bS��}�t>I{0O�D����V����Ό�5�|\��lχ���Z�DG�@��}��c�����ƻ&s��?{��p�{/�lZ)���b?!�غQ�@�{��)�X�-�\>2	k1L�x�		~��t[��d��Rtj!@�o5�0TWm�X��|����KBs��9�9�̚�f{��und@%���$�&���lɳ}�k=]Oӊ�N����Pe+���KE�����W]�@?b�	�d<�+ɡ�-YF`�����4�:���X�<H#�x�E �)�?Ӄ���rJ�=���zI(��{q�2;���*� ,p+��ة���uoB� c�kL�J�Bp;O~��Zp4kt/�?4��7/�El�Ml�&�j�rS^��?�S�|O0�1C4׸�63p������s,���%ӽ\��·��Me���� ȫm��[c2�gx�G��_�CCaY������<A�����5�25��x�\E��W'˧􎼞*g���Λe2E��D��v�x���4�B�R���d�jm��q;~�����K���dV*np�E��D�kWXL/�b9�+��X9�����m�p�E���ɘ�-"��󑒟�8�����)p+����\�;+�;�⹠Lo����5��u�W�#�q-� ����W����X�5�_�D�M�۳}���t|v$�*�唼e2�XgŽ��ŗ�p-1ea�i�D���B_��}��$ƿ:��I��Lt�w�&�֒�(}�e��H��r�&��.��d����\I�����)�v�����8���l��-��F�|����G�/Iay6�
HaP67䂡��{�� c!Z��\Fd��\[w�vj��"H�WrE��V&��6�߃3M���R�U���S���0lǬf�kI]����]�v������=��	����h���f��L�Y���I�T`o���Tl�J�4t��IƏJ|Q��nmu;p=��)<�����Y��}�u��[���� �����^{���]��at{�<{� �F?:�@`��K�vH���y6�|����
9�ݭ�Z�s?�m�ϣ2��!A�h���F>��J��R ��e����j�|���\�m�֜�DУ��8�0U_~��4�����A���|(<�_�؎��
4���C�XE��l�3�	��(6Xj�{�n�>�6�@E��4�%��{s�{��["�����Xy���&�~��uH7�fvՔ���wkǱШ �ߢ|)q��;�&�YD�T�ĕ�5�7g`��=�[����ق�U�#躹�4C�K���Z���J3ܘGa�/��,\�5�2�
�5@*��L�����J��p�����H�ցj?�eAFi�H�����*-��k	X�ht|a���z�#_��o'�{���ؕz~�8B�׉�:��&�~�d��2�^����ULp�0��Ma���̋��t�̵�J���Z*E%��~�\�I����;�ێT(�)�,~�N� ��Ց[��.�+�@�Ak�ƽ��-��>r�Ij	Lr��o�˶�� ��F��WS����[�,�2~Ö��մ��&IM�	�J�M�I��SB-b�r��o~�s�x��F{U�hV^������>^!h2��d���@�SQ~˹@3�+1,/���
��~C�q0�~���z͆y���G�j�@�Y��e����i`3st������.x��;����YP	\JYO���w���~@ҟ�K��4gJ�;�t�g�ү�gHu�zV#�d��S��_� ��q(�@+-_�hL�a�Ln?8����U�Ѣ�Zᥪ�@Y�֔�NV�O!���f�UA�p|Me���R@���m�J�]F��_\g�ha�̫ċm5Q��e�mE��3�$�t�����%�S��Y��ƒ�����LP�R��P�!:d[
/+��B�kX�R_��ZB.W©�!1$)�J�fц=p7�Ҋ@J��S������/�<8t׍q��fj�㔄�Yq�& %�7��W8$��͙",�YG6��L(ʛȫ0i���C3,"=��mN���p�Z1�o�"�u<>��w9���e>��J��T��"��@V���=rn���E2���q�Ƙ�dz�Yr!I�%-嚘����~���yző��#7�Hsj�d.ߚ��������U�J`I:ן�T�%;���&>�����૯݋��N�/�Җ(1���7$�b<YM�s�wB�E��3���F��#��Ģ�epWMø�X;i3Io���99��&��UW��wO��g�͖��֛~��������a�/\>�A���>�^��a	�;Kh�t��Vc�4�[�A~���@��S��{;g�Đ
`̔�{e�M@y1P5Gh�4�� ��b�+�D��=ܰ�Sx��t:��z�p	�!�Pa����H�[jC0;�×����O���Qءl�G�in8�v 6��}Η���+R�D$�p�����8v��jX�5e�qw���Y�Ϻ����0�����X`�����Q��t�^���=��ܷSA���*�^�`UĒA�B^{q2�Xd���]��jrHO}�=�ZT�b��e@U��M�&�+�Q�c��B#W���
��%N�����#�-������T��Ǥ���;Ӆzƹj	p�u�ǵ��?��L�,�+�7QX�/�쎨�1$J+G���+;c� �K���
9ւ�P�9(���}Ŀ��J)��[�C�y�h{��>�!�Y���g��d��l �])EJ`
q������5@�S�ri�_���_R(;0h�:[ �Um��õ�e�q7���W��RO��{v���/q��G� S�țl��Я洌InÌ�I%c˒>Ŷv�P2V�,?�K;�K$]8��(!�r��%�2��p���}�1\�,��D.�9��fw��u%U�y��hGޙ���12'J:�Y�}s�� B��1bƦ��#�DJ�*�IO�-�U���=�3X7!��<rAe��f���֥Q/�c]�(�����@���pN�c�_�d��������� bߔt�@o�i���SeH��ITJ@,�q$�b1�W3�ҟ���g���m��:�C幃�ŵ݉�����Y*1{�]���\�����`n}9U��}��CE�Q!�OYiU/s��%����N����5G�yB�haK�oE� }���㔅�!��NF,RJ��I�Yѷ&5*,�hI@J�+�e�l:��{�ص�MpB<Q�H���5�y��OJd��
��yj�`4ږ�����J'�,v�������.�����h3�ө�"/��W�Jt�"���\��N&���<3�}��n�ش6�WCp�e���ۥ6�{��P=��eeۍ�}kx�ڎ�����
�Ԓ�?�K[��e�?^�d�u&33���U�Y�qRH.�W3�2�4П��ɖV�����q�����b6�5�FXx�O2��t>mZq%���'����nD�(&���z���Q�cb�zn�F�L��w�U�^��8e�ߌO�q͎�j�٫<V���y�V�[<"�'�jzY�"�h�g�`δ&9�s�!(E]��{G��b���x��!4-#Z���w�v���˅)Ĝ�|�g��$���l���S'� E`��b�+��N��d;BF�"��&��n�yz��bc�wB9�D����9%���憑��۝��w��8��b�&㤌g\Qmx����N͕;.ҋ�h�vd��1h}J;���N�:�	Ed��&u]�VVؗ������׮�!�߹�-�r[y��k���fJ����l#�eo_k�f��ʻ��b���5F���~�ٱ��Z�h��M̾�U��:�&>��1Ld�\��9w�с�)��t"ۗ.�NSpP��bz�"X�'����29�<���)_