XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����#�5[U�q�# �u�0S&�r���b��řI�Od6I|�'��	�BL З�[8t����{���n�el��sa�xD�:<ͫ�2�x���:�g���A �:X"��5��ɫYw��ׂ�	DsK�(/�H�}I��G���42��gW���V1wd�fS�,8W�A�r�D�~���4ԧ��c��[��#?j�A�e�!|��y�n�7A�F�� ޻)�B���T3=�21�n_Z�~��4��J~� m�0��v@�����yo {9���XS����~�uV�����gwu��a9�\�?�]W��{�!�)Vz��@��]E>����R���"v�ؚn�e�.N��<
���§�~�h��Cg2���n2ܺ;���[��9���
x��ȅ���n���kT.���;�0�u��3�zZ�_�y�V	nl7�lV�Y����[��H�`�"|2��a%C������4o�����d=�1Sx�p]k��<�U�_�Z4�4���7���n-2&�P�J$�|�t���i�� �����4�8pW�U��v`���W�_���u���l�M֔b.�8�*]b��>>�D�x-V��fĢ�5r��p��}l��%0`E����������9
��Eڄ���xn[ղJpL"z2� �a��S��g�r�oMx�9�����H��l#m e�r����]��,��p�i�� Ck���rEa��%a ��������)z����r�v��ӯ�C��{P���XlxVHYEB    3da6     fb0��=�L���x�ڷۧY"a1�s���q�9�PAz?���`fK���׉�m�|?����Z?_.ְ2t���� [�[�A�/�l��ed�|��< L�f$��=)B��ɺ�>���2ͥ��KW�:�Pa��9떁&��&{�u��Ӝ<!�[*kl���Q�kj:���	���Vn��E�r����k����n�����;(G�T����q1����qbs�(+�9���nS�֬�H�!���$W_�r!b��ٓ���r;�}bjNr����ٯ|�p8��H�T�戣�6���B̔U8Q�1�F��8"W�BX@���E�0͔%F��qXg��J��K���'�� ��ҳ�^as��.�T۹�xk�J}�-#�B�q�S0Φ�E3������i@�spY�3�ރ�֬K��"��<�' ��JHD?�#�CYj�x�s�ӿ�[��,�Y}p�F{�;j-�R�v$��7�_�Wh���۬��1H������a��NMN��ru8/��(�8���z�7�9�X�VYݜ�NpFz�m���Em��L�ϰ��:�Cx�]>�!8[<| ��aR��GƄe�r��w��%��P���5`OĖB�����V�5ϼm�����~ec����XV����<�;�BDW�*��r�=Q�Ζ0 ��^��ZϏ�m
5n�O,�J�p�Xe��Y�4��+�%�>�Vl�n�������_�}8��BG�ڋh!�v�v�":0èj%o��f�T\�-�g����?o�hQQI��}��a���>A ?|���"P�n����8 ��0��
'DM{b�|�u���Z�h�R!����O*�Z�_spW>����rR�ձ�C�xĲ������9��&E6���3�K��L�*��!;�uS����`�����PQ_ �$G+� V*;{,1l���t4����<��8�f��pP��{�:�Xkic����]�"��ׯi��YYX04ə���;8!if�N��*G�/!i0�*a���қ�_G��j�V��(S��M��s
< ���������!�K�B�,MO
۳������`��-t@�s�
89�j�Û��EEü�͌ ���,Q;ǭ��*�h�{^� �!8?Bbh���ΏX
�����_�O7:������R	���DM��Wdb��r�
��ʇ)_2�جi/�3g�?5��Oo��ΝC���jЀ*Z��o{w���l�h�h�Oc^^�"o��UN7�/��%���s@S�)�3�0�I&Bə(�[�4'���~��u$�8$�$#��k<��t�B�e׌��4Cn�z��E�{��,@L6قJ�1��X���<Y�g���c�56վ-cyEmԅ�'I1f�b��x�&�{�%l�yN�۩-�Ɍ$~�s�������E	W�x�d^\|���on�`�hH� L�Vw\`!�b07����",�=1Z|�yǵ�ܒ� �2zR^5��#�JQ��8���WHish%��y��:d�hQ�K�A�a֖#w��L�qV���Ve�V�X�=!N�HEG��`�@Ő�H�e�K34������^��Ug��j�iI(`Z�Zܫ��y%��6�!��S�v�!���}DE�4L�bA}�����oe��~v�2!��,�i? q0v� ��!`<<��nb�xd�<[�Z@�Y�����[�\!��V܎�%���ͅA�ޑ��̢W�_�yJO�{������A ����Q�zόV���~E�����!�jb�|΢`�M�ؔ�	���n����׌_��u�h�_f��w��d�����^��{#���h~?����y��6��)E_	�>D�/��e�r�U5�T-���9�#pkFu����,Cɟ[1��\����0b�W5n�y2f��s�z���ѹݦ�쉾.r��o���
PL�b�h��ZX&��u�H��=7�{&W���I��4��S� ??�����z�����{!�o��MJ�h����cZ�6��V�ŇTD�ؤ+qoi�K�&5��g�?7Nﳂt��	��D\��ॏ��ia�0��AϏ���E'2m1�#?��T݉�d����(�T��k�i�b�#|�3�ۤ�h���DB[��A+q�FyYo�K��,�j*JeKUD}^/&c[���恦��.�_:j�H�PQM7����$:�V(i*�diq������@��AW�_��u	\���� H��o|1��=n*a�����	�
�By�[�3q6��X�kY�[�F��l}ّ��wc2]�H������(�˼�b�3�֕)c�½��/��<��~��.S���J,����@�F�����C4���8�����0���P�^��30��lLȔ3�ń�ƽ��DzWr꽉s���&��o[��~��%
��o��/�tUC��Kd��SC&q��R�� r�*>Τ������әpYq��*��0�6j�/ձ���6��̺��<�^�,�����,͊_$��yQ���j�(m=������3(��&c2��:�L�t���iܪ	�+�<�[,��~@Y�%!�����3]$�=z�v���q7��>j"+�Yq�$���LCS�q2[�1�h�ː\:B��öϣ��<���Y" ��\�,�@f��nچ[��BOR��N�y����� ���j���@H�(�9u\�>F2����d�}��7�i"�[���W��Ԩe'�Ӊ`-.�O\Ƣ?f����6��E�$!l��5�$�2��yJ4�DVv���](�.e�������v
�ϨLPƿ��f����8��~ߝ�CPӅ���S@��;�#��X�ʔ�X�j1�]w5��q�G<��5G��{���������r��^޾.2*�=�`��ل�?�����ִ������=ڝx8SëX��\��U��@�<}ye�h���A����kNL�5S\r0��x!��&����yCL�!�QA���O��4r����A%�c�[y�˭��2��0IӇO��Β��S|��ڬ���Q��=��?4�"��u�c8�˙Ip�.N�1E*�@!�$�_Ԯ�z���^�{+�3 r�����
`�B)s�����Q�lC���=�G�.�O���AZ�>� r��1��1�%�es��9L��9 ��j���J7q��ܐ�O$��X~�Tj�}����Y4�p�)2�S"0LL�C��`=�&��k|*gw(��<�%��`����`K�Vb��8O�A�1�!vy$D	��Y;xC��-� 7h[���W��ѐ4���2qv_QȗC�1Zg�LT�`6U��p1����e�:��o2P��q�d9����d�L�����&���z��2ړ�P㨩���	��=2`^A�}"��H#��A�:�hq�z36�`*F7��}��Oz&]�A��E�F8�\'���HA ÈP���"��2���Mn�E�8�'s�1�^����E2���p@�j���$��y|%[��~�f�N��ad��]��5Y�Բ��k�)��������܊�u'�W��ϣ��r~,["��l��@��7.�&r; 	�86�Fe�F�k���hnZ�!1k�3*�3@��n���;)��%+X`�|V�1]�eX��n?�oO�m�t�
���F���2�������]�2��_��ܧ~�CIٖJ�;��,Z�-�ݐ��0�א��p�s*?o��<�~s�q'��+���ի�]P����µA�R��mn���%�4ƻ�οuSCoY�>�ݮ���)>S��7�B%&��rs�]@d����xE�ٰ ,W�"�vd��ěȫ�dg��&' 8�dQ��a�(����L��Agq��̱8�e)𞶍O�=�9ֽJE5J� n���u������G_4�9F�|e��ؽ��S��F` E,G�6G��c�/��<:�[����_�9�Ϥ7����ݴLD��Z���4ݮ����Fa˪���9�O���Iz�V�w��OE$	ϴ��u��V�$���1���1r�