XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���;O���ՙ-��+�E�N_�l����E{�(���o��q���כ	6s��ϐ_�c���,�Y�����ю�Trh���n{HODa�u#��j0�W��g������J�H����I��*��\�t�����gVl|Zw�mP�c�謆2fp?Hq�;��896JVs����@�
�L&t��E�]�h.�a�ʚ8�y�%`�׿�l/z�� ?�K��=tv0:Ъ��gl��\8����O�T o�[*J�f�X Z�_h�
��B�tR�8��b��6�r����^����&����=�¸��Rh�̄�3�z];��Q>5zˎ��n��g��,�x�X��P���Q.@�$Gɖ�h�� >��Q���KH�wj�y���I������ж>l3�����J�Fmv��OW�z�o����vr:Z��Ʋ�8� ϡ��X:���Dt-P�+>�nn`���t@�Tj_�qB[��BQ��I�k��.Ǟm?� �'��'g����~p�|��&e�f�Æ<_�'�W��RJ�΃�{o
����#`�����ax��eM��W��H���~���"�(`8J�Il֚+%a�{��+��e9��"h�/S��!�������)��gT�4�_\Q�q�����RP���j	���~ �Y3�s|�
MUW������.��p�%�+��Ld���WuBC�FHڕ��9)MW��q�a�	M����xȁR���(b�8X�c�1����}	T=dU�XlxVHYEB    dd8f    2160{���z6��Z��kwS�і�L�����K_���Ŭ��f�>��@��ml������� �q�=!rg������s@��mL�m_[��!�R�;��ȉO_�tu��H~�k*t�o�x@�&Ēt �ü��'!�O�I�7$�����0}K1��۟F2�V�Sk�u=Z�Qq�>�(.0N���B�]��]�h;- jhi�r�f��.���M3݁m�ė�����u�]��$��a���X�eޥ��l߇{���?=��%����́��>�����Q�U3��"�Y�P�9!}���d�3������9ݶѨ�s��yIS^��ǧ�qn��op�k2��|C�� �%ZN�tqC&�P�RYRa�ٖ#���c�S�mcAQ!��E�̂�.�}�3:�q����"���T�P����e��!fǓ�k7�n� ��A�Sտ�+C?�-�Dj�L�5)��7�o�(<=�	�5|�W����X3�;w~[���RQ�����7T6[{P��Ō�\���l�[�k�0Vg�
�Q���%=�<�8�,��4�g��_�����a��$$�|P����DīR�"BV�L�ɕ�%��ͅ ;����R�,t�9r��(-����m�|�{I��y�ɘ�L��G���4Q�Igh��A}�A���-��A��O m�e�Ъ�^��l�����K��ֳb-�����z��ul�a���DT�FK�Q�;��F��;�[�XF�<�a��iJ�����u���t2q�_Y�3��%�����2�
���J7����o���3(G1�^>��}��6_ߎr-����0���:�=��?4x桟	� ��z*�B�ݎ%��T,��;�gG)a2Ǝ�s-���GV+�N݉ODz���4	o�黦 ����J��z�y��)�!�ɂ%9}S��S�� V���a�p��X�^�g��������LV�*b?3�<^q�k*R��OOb��0w�MZ�qw�$�׉����y�m��ab"K�@��������^E��Q�����_ym8)�!�ݠJ �ԥ��m'��)��E'����;Y��

e�g�����k���m�"[\Z�[�{�;�7{�h��ڑ\��?!�m%��#'�s$��;U�Zd�u�.�J�I���u��R�&��@o$ὠi0��'Β�4Z�B���c��<<����m2�#�c��"��4�2
˗Խ`0*�ia�� BK�ɍ���9t���0E��g�Y����}��*�dQ#�l�����?��dS�2�}v����P�����9���}�g�{�3"*�_#C�ӷ~58�ܰ�X=K��� 浆��k�	����#h�KVPG�<����pL����
Z����ܦ���G|���
��^� ���s�PUC�[��������Pu�>A*[M�#(1Ĝ�P���G��4�J��X{�l��$K�-e�� �K!�s�eK��/U߁�m@}����$�
��$񃩏����P�r� �}ʁ�M>f����H'zt�σb�=��쎵-myd=u�JexI��@� DcX��V��ދ.�I4l ن�Q㋄P1���V�����L����u٘?��_�|���U�1�Ak�д�/|��G��lo񎁀$����{�����c
s+��X�V���Zh�i��'����G�M�Ǉ�w�k�M��.j�ۇ� ��7���7�WٶT}�n����]t G4AI8K� fN� ��t��$�g�y�n<�Wn�A�2
�k=_&�J�!2��,�DɄ�:�P�$�H-���W�B�Þ�n�,�x\�v���5��Ѣg�ɊxGpE�";ѳ��\y󽭝����eby(V�`d|�(�hde%H� T���R��Ks����J��mh���c4����M��ڝ��#_��] ���^�:ݵY��.Va��N��MJ��A�0���s����8�<Ȝ�>5U�uJ�]�R(D9� %uG�ܻ�-�q;n�ZY��C)ao��I�v��>�rb%�pv��d�-߆驸m��9�FU"oh�|p=z
n��!��<�ʍ����|Ra��*�>/�[�P2�RR<�З��%��5���0�Tv"�l? v�~���}�S+I@����R��H�RT{�6��ׁ���r� �e�J���yp'�������.X+�	E/N�r�;����g�
Np�s��)/��Z�"���jנh�"c��o�$P�a]ߊ�@��-���������훈�O����dl�$�)��ß��fD����ʥeE���u:܉3�<Y������Ĳ�� l�7����g�,��j�mh��5��)~ ��pgʄs�rb�_��J��V��X���x6١r��˭���yl|�Dt�A�(�\�(�WP����!�W���UBWL���F�PNZ�; �7�ؽ��������ǻǡ�T�a㋉�U
���w:�1�ae�,LW�����(C����ق���_��j[A�+��5[�l�mzKS�12��O#")�Y�;�<� +z1q�XXP�w���a67�߇��+V��\Q������#�5�X�+�bZ�T���c�cǡ�����GX���$by�ab��ݔ#	N��AȌ��'B��t��U���2�ʚ�gq�������)����4�ꆐb&�f�!���6e�{CJM��FDa-X��ĉo�rQH�R��8'nCg.�i ��/�b�	Q$��E0J���2��}!���>�T��&����f-�RHEM{�cU(�@��Z���AB?�P�`��m��!N��7@x��4�S��DsI�=�/�!p�~/-�����ң�����yb���h�S�hY%��Aʵ�׵�V��w�5�� "1xi�+;Ȉ��2��<���:��r<��s/�^Y'�)���'3W}7�O�")�M�tČ�}ö�~IKU�W�C'l������ɂ8��5 �d�
��|����c
�uc�����ReC�F���QWÊ�8O)�)�`��m2��s�=#���݇���!R��9c!��-q<6e8t,�x��]q���o%�y�YR.��<G��?��l����f@ܜ}���$Ƽ�\�K��
�d8<JU�q&�&��K�j��;��,��2�z?<��CZƌ�oR�4�+��x0�Ժ�p�[�gD���Y�qOեg��
,Cd����t@�^�Jh��R�	)�q��>��~����y-�4�\���� ��K M��U�I��py3¾_:1��$���Qqj9�����%%��t����<�4C����p������~Vp�[K>觞Y������V��ӳ|7���@V�+؟ʆ��Oש֌�f1y��@�>�4��+,S�T��K�H{{xg,	�gkӥ44`/cKC�6sc�-�?}�A���YiQvc����V+<M�*�HL"� ��m��b�`Z!2~.�BFQZ�;O*rDc���-�%B�֖D��ycb�P����H�$�b4PB�CZ2���o��ٛ4p������.��\�N�e?�W�Fh���S�U8�]�]�އ8~9ސ��԰�F�ǿq#�I\l�̲�{_�l�8.+���C/�Ł�<�Z{�.^.�̦U7i8�_^/3�v�uj [�`hr7L�a�j�
rS�y��7�� �tn��������o9�w՝?����F�.�vޑ3��Г@��J#�}�d��I#�K����8-��:�5d!�=j� ߊ�%,��r�p[��#V&Z�9�����e"5%'{�U��2�l����^��Q�K9�Jt�F�׭i
8VQ�>)���Rz��Ŀ��܄�a�<�P��(������Kn��F�������{u�ٺ�u��%� �,ʊ�+�2��-�B�q�ﰥҝ�V�hnW��;Q�J���a�<c����>��3^u ����6�Go���RH��({���3�u]!Ye����{��)�k�^�v:�^�����9s��q�����тywi�v6�X��on���Gw�H�HX���B�*�:�5xmȏ��`"��;\� �G��o�v���)��8��)��*�4�f$�w��;Q������������Ux�-��[%
��J��3_�X���S��Fn��8������E5�((ʣ z��N���S²/d�?A��8ĆyBY��%��g3P�q�#]D#��i��.����ћ������5I���[�t�?mѵ	����l�Lp̛K�Swؾ�p�Ȅ��8��⤉�c����6MJ�!�3��K���U�� ���lB�h����$�`V�9{죎�9�jv�MV�!�O�2�����H�Ƕ5)7���!bqjW*S3L��U]A�8�hS�3n��Ƃ�����j6��!�ci��\���h�\'�R;�M���%�dd2��W;fd��F/���5���E��HO���U[��I�H�Z�fX�6����\0n���|�?y�ϰ��E`�O!=�.m5�b�!V����� �C<��!���k�ѷ�n5b�bv���I��|�]��W�ڵL�$�6�|`�v�	F�V�w	�
K���[CW��0�^�Ѹ��7'V#�7���L�dBJ�G
��P��ޭ:�-��^4��dmv�TkI���	�@��9w�Γ�`{?��j�;
!*�V�A�,�t�9]f ���B��

O���h��Mw9��d����������A*�{��F$��FB[����Ħ��*�H��n����W�8����Y"Ӹ�M���ǗS�G�(���^$
p}-J>�8�r�0*Ypߐ �;&k5h\�['/�������-4�{�H/8�&��ޓ�aI� ��̃V���:�Y����X����(!Q�O�;8(��3�q��]�X�>��ZpQ�,D=j-���zsV�@�����*�����(�O�]˃�����U�r ����?^�ܛf,�I9F7�\{��=vCَ�0��r�/���a�lq��p4��z҉_���Y�FU���Wt��V�Z_��=�W�nդ�ܑ��n��i�Y8Sk'��R�M̎W����g$�̕�g�Y���(nCm�(8� ��u�j�Tm_~�|�j���wN^T�wF� ��N��'ߖ3�ن�A���NN��T9�]I���������73���Pl�{��A�`�������Z3'���Xf��z����6P������A�̪���m���!肮2��>�M����ݪ��89H��4��wqv�vM!h7<I᷁�n�;��Y҂��
*���@�⻤�W�Ε:X^��aEXk���ǡ��R�]��ѥd�b�I%�UI���.���S��8��t�Z/f6T -��bT��4�6c�q�Ħ4f�Y�V�O' �*g���R��ʒ$����Nt�����Q���Q]�;;D��@�{{�~�K��Q偏򚚸K=��:<֊Χ:G��xp����l�ŗ+���Dr����K�&m�!��J5����,��D'/UdA������$q�R�P�z|�X���@�4Z� P�s�lё�vk]�%����!�=z�3�+?���bڷ4n���|(�ׄ�9s6��ʰ��h�HM��3J���z.>�/�4I�KE'b|i�dk�����!�I������![�@o��m[�k��&��N�����T�=�t�A�������I	�ySg���|br�2��*���lU*@�V\)�'C,"�znr��)��$k��g�%]$m�{���b%r�sD���P@�o��RE�5��-F�V'g?PnO���p�4�L����u Jr5�H�ؕfS�|`HZ��[�jj-������wt?� ���m�K���/��\�m�@�jت���5vr`݀����h��a��ǋ��BIZ
=�=ɒ�aݢ4U��K�,�y�W��jj ����!%�	SF�Xc�ӎda��(6�10K`�>��c��?��@������r��k嘋6{k�_����
7�9�#SV!V?��J�3ar� ��h��`SI�g׻��$����GF����[�K��PY𔒅���Uǲ���iK�'y�B,�y�a1���#o����F2��v1F3g{�PJ�X��iWER�@&��x'̃x��=����cG,��XdX�։�I�^-��/�%d+q@wܜ�g9"�ޙ�m�*`�x''\;��#��xQ?�ΨJ�Aͤ{���2b��c�B��V��)���W��a���#�FVn��x�2` �(�[��=Ϝ����Ed�J�~cx����l����`.��4���IP������r���~rzæ5���@i��Շ�������_��}���#sW��ټ�w5[䱣r�����ET�s�}�
n��W�g���\0�bW���i#�b���mɴ�9Ji�������*$��n�/Q���5��T�`��$h�T�[$߿�^ ��_KC�W����s���ѯC�QI�r4�&T��b�� �Pe�c�֮U��8��Gv�>h���
{��{)��m��FUDc8�a6w��{���+��/n���x2�qæ�lHk��@�X �⾘��J���-�f�s ��]1(���}���6�p^�enN�ȏ��������1Q=i)#���~B*�G�'&��f���M���f��u� �"��6��^O�Jz���Dʙ@g��2��.�f'�͌%g�t��T[2NQg�<H� |���+�u��i��3��M֋r�L�/ԧ%l\���4�)��p���Bj�MxOMF�.�w�����Uz<|��eB�%<�7t�ٹ7�?2�߽I��V�GQ�"X�}��ˁ�,�����ĸ�;<��ߨP��͆�V�[�o7G ����e8��CWX[����y[�~͌�;H�O�e��z~ ^��ْܣ�>z��3tLAޘ[�B^L�R�+
wg�U�wC�%���VK�٣�6�;=���Op{]AyXqQv� ���w;������]�X�z���rv�@�Nm�NZ5�&��2Qt^�4�R�:��=�(���R�1-�M[e�KN#��9�:?����:;@D��l�F/ޢ'�S ڮ��g�Kқ����zRe���=^"p��?狸�M?aJ���y�a��i��K��K��o+d�1b�G�j_�C��v/�`�n�%�c��ͯ\E	.	��y$k��X��i4d�ᡩ�ohR諡8�q�Ā��J�%���������)��ٯ�^6��J������.)��F��3*�ڽY��cY��7�����X�ʼ��s�td���vES{�R*�p©(��˥��?}�`.&�en7K������ +����s��/*�A*��I
��d�BB�*��Εk� a�k�6(��gM�-+�5�ނ��,�O0���JQgU	o4'>��ږ�Ev�s_��j3�C�"cA���8�_Sv��ߌ�Y��6j�/w7�r���IQ:;d�I�x�$,�9R�s�(y�VN~;k`��Cr�ah�2���N�
��'V���^� ݇ �C+R��g�z��M����L���شv��H���.��Qm�+���%X��X k���w�����3��+h���k�x�b�v4���іQ�a2�.�g��[���4�b��1���]g�p(Ʉ#ߌ��7b�na�vۯ�ުf���N�(Φ��㺵��P^b�� ��I��=�^���tT���i@����<�i*,���!9/v�c;C�OM��8n�^�L�P|.�&<�8�J�L���O��6�1Ƹ�J�l����6t4��D���c��av�vt�0������ۛ���^!:��+c�Ș�G_!���vA��L�؝f�6C_g����|��<ڹ��
w�.	�v�V߀$�`G��r�.x�n��
{�YB��Oa�音aN|��ES�]�����a��rY��Bh���J##�y�N��HwќBJf�F�ڵ��JRtk��$�������7���	�� ��}��7~�H��E�k_#�/��/�ʾ}Z�	��&��h�2,�)�����&��Fβ��Cr-2�\F���q���bh��YrZ���ҜS����N�H��T�D��t=,Q����gxc��j�lh���yఠ�F��/�����^�Ď�l}��e�Q����V6/C�����-����#��#[��h%b�|��r�(k?*Q��	��y1Y�@���k�����;p]N9N�p�N������d�PMI�j;2�!�"�^���d�lz������=к63$5~�U�'1[�j���M����QTl�S[I1Qv�}��#6ٮ�(�>T��`�sC�@���
��=��c(�.Q�x�b]@� ���a !l�F'G�#.d�Ky��=�Ϯ����og��B<��8��3�["�H
���R)j��,���H�$l̂���Y9AնV5�O��0t]m�L���йb3Kr