XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t;T�� �C�� ʄ�1׃z&��;�|� I�p�F-�y����7v�X������螥�#y�_�\}s�� z��q0��C5*�d3L�\���wr!�#�*���-`S :��
�S2#ZK��B��r�f")$U^���	�}���`3Z4��D�Q���!D��	c�j��q����Z����Xa�f%�u�J
>,EN��-V�]��[�w��$�:�p��'���W���oF"�
%���}5��p���%T�T��"m���k�ʆ����G��b�N_i�8�K�b�a���D�=ST2�t�F�ԏ�U�+�s�ʄ(JM�],��P��P��Wg{Aw�����2Ub5�����L���癔��x����	���?��j��	Ua�F		�z����h�v�P��y�a.��R@�s����O�kP2T�zsؕ�Q٩4���4�s���~�竁�7�X$�!�;�.����gS���`������^��p���M���V����DF�Y��_��`cG=���q4��ȸmk$���~�J<��:6$<�{��ԝ<�Nu����39�+�zw!�|��u��@$~G�
�j@|R�'��B�Թ��6u$��;Vr<(��M*�V��+*]����:�{z��KxU'-3Fw��ts�H�tJ�
��1�e�����+6+cr����-yݰ�J��sU�$��(_��wԝ�m��*��Aeӯ�Zo�� �-���	]&_�}p�T���?=O��$�%���XlxVHYEB    b087    2540f��:��]3{��8{���O]5٠ơ�3����4� \�E{��AR�;+n�D�r9 )�3��M��ab� �O��'���VER"t���M�	B�3��q�@�������i����"�U�����ߩ�b�p~�3x��� �m��@A���:����ei�*i���:����d����h��v��~��sCAI�fQ�b�~�P�R��O��O	d&/�z�mS$��|հ���R��{�\4�ƨ:{�����{�c3����!�Z�E�P���^Zjv�%�"�_lz�u��2P*�c�z���۠�s{A$��7���;m�[d�1��:{s}��|�r9���[{,�Y86_7t�i�����!G��q���Iw��g�*S�Np���W�㧦4�(����ʼ�u*��uC�&�}Y����' �G��G�:�Pf�=��(��M���3�/�wo~K��I��#�i�d_��y����X뫞�_ȋ��Ȁ~OY:����=X�4M� ����.��จJ����z�?.
?���S��@��A�Kr���*�5z�ã� �Y3駘�?�o��0��Sy�'����<��t�?��K���=�rf���u+�;�2a����G�R�c]k2���MC��ϙ3�q_+xmLh�������r�21��W��ޙ�DV���+fн�X6�v�{�������{0�sFH��(Iԩ�H08�4��^9N/� ��a���N;}��`z�֬�A�T�K�\G[Z�2'��Xp4��,���T��s ���aNO�#��-������Ġ��`��3���\�O�A�O1��B���@�ne9ݞ?4�N5�>���0z\hZc��a��z.�?����d�O�X���3=��D4Cr7ܧ�<m,{��Y��5���zs��|���ޞ>����[\�Br�
�z���2b���h��d�9R���Hނ����u� ��8s+o��'+���7��	��>��P���u�M��f����x�8�0� ��)O3��Tr��&�����y�s�_Z$��+�ȿ��`ƫ���UX�b6w3�͐Q����n��_f�ى�����_�2���1ϓj_вGo��7��-9d4�p	����H�q��S`��m�~�^�I���"x�c�7��ﰊ�sc��E�]M���w��])�"MS�UAw,�6
Gѧ (��A����(<Y(�u�3g���4���z�sULڙ����r!�xk���/l������(�p���<d;���i݃gL��˧�>�]p>}�5�Ǣ� ��1���\|�s|�e����@E�E�E��R������r���?��f�.�P�6�����1O�p �7��$X��!���3}E=����^*o,��l��j��F刷�T,���㻔N�˲�5vGvH����Zх��'������}��ZM��F���H�5��Yr9���i:��ºKZ~ɱT��ʌo�+�R��`T�0+��¤�!���W�#�M�y.	Q��hyxX�AF�ϩX�_`G�eeI���
H��l����@��F��;�Ͳv����m�|c��h�?���彃L�eg��>�S���+д��B�$���fes��7����S8;���d���c!�~�B�]�S�$��t�N+Y�	Y��a�Nt���@5t���>�#E�D��` GҊ(�ٞά�8ֺ�Y�[M�mk-m�~g W�3�=�j�֤���V-$�ҵ~����t�N4��s}�>R[,f����y��L�u�q�J�j
�j����9�*���r�g5%��s��'��g:A~mq�,AV��>�fm�l�t��^�����s� �Vg�YG���N�!U^�ԁq!�i�"��6t��Њ��CR!�0Gk���O�'`G�@���&c��]��.^ܧ��^Q��!��:��7�^׃�6����γe�c��Yl\�|��W�J�g����!�� �5�Xw R�]����xJ�$�.��8Vh(�,~���h��b���N������n���!U�3=�"5���U�m�������zf�·�̝�ɿfX%`�+_�_�_�yt�.:�N��k�B&W�+S�|y$��I�4q��_���DL@�z�-�ٯ8����Þ�&��\��H�<�C���<��ȡ� d���B���],�
0B��D�"�I]틤�<��Ɣ��Pfɯ|� ��k�;A��i�9�Rh��4���ww�:[D����®���#��������<�+'�����<�.��3�ʚ����y`���e�cT��a-+�6ۃ�W���c�P�x��ω�.���6�T�7���*w��<i5��˞k3��cWL;���:n��zA�.�N��J�ù5�Ñ�@�G�ܪ�]M�U�Ы,
(���w���}Y:���������A1ܳ_�B
|g
��-����|.�9�)J�7Ч����^���#�J#�_CoxR�H�4B�t�t�AM\���g:�����k�D�x��.�
��v�ՙ���(���My���˷Fj�����]���ER�\0�ϜﮂN��Β��)+NE*�(A{��� lV����5���4o%i����;rҬfs��]�!�x��L��)<K8fM�(�u{'��	��I���7>������_�fL~��^/�2^6�K��o�],f�O�Q%�?��E�^��� *K�՘�$�b�8ƈÂ��Rn� �(��m�c���}�yp�/(��>6���� JQi���_I�JQ�iF\Z����)�Z��qQ^Z�c���Ӑ7�܃���=�3�|�5��~����|��1��Pm��t��߳�_�Rw��` ��X�L�E�t�2@���D��Hc��S+��?E�\!"��Po��Z#�@y�?

���'B����dt��=^�
(�m5�u���{���]��z�0�s�y|�
2����;��5��j�H0��ה���S��=�l)�J��r7�M�f=���H����+�.���e#:��lU�P|�������X�b8;I�ld�K�[����`�:�9^�6_���6I,3G�G@���9p~��~�HV�oϭ.�`@�/>�-D�hW��c���! Rё�W]6C�(qYa#��yd� �٤�lhk�y�µ�,V�IA%y�����4l������-a'��iH�l1^�>I$�u�i��)��T)A�K���E���'����b2���{��L��B��~y��sh��r� ����yYqno'u�KGT�tB�� >��>��Y���D��ѝ�t4���5[+w���+�D�Ok��<cKAsؖܚ$���s���M!��G���i�h���%ְ��>�9;ao��4���F��M�ܷ��
B�Va����Z�k%gʤ�v�~����9����6��­o3���H��8�@�MY,Hɀ��r(��0��Y�R��;��ن�n���J�{A�5u<JO���E\��,J��%��m��t	)+j"�.oӇ��(;@������Ʉ7�����QQo]+j�!H�'[�p
��.�l��>��`��}0G �� z��ca_l��um0�=T�TbV�ΨnycG[J��@1J�,�����qZ
E�|&������:�� �����)���B�k��T�-k�(h�ҕk���;NX�;M��������T@7�("��������I�b
�x�@���w �$��|����4	Y��Ɩ�-h0h wUh=>t��D�{���b����}��-JCcǧ3��NG�g]�Q��4�{���uT��#D�A8M��%U�^��K�����@�F��R�g�f=�ty���|�rb�I�;j�����!*��.ϵ���B��(=v�>\��[)e�/UЩ�o��v������Z�b�۱��F�������1���Ӽ��z��$4^��D�` � nR6g���Y�C��z>����3�<(ۣ����
Z	�?�@ބ]}�xB��M����%7&�)�dE[���/��٠;"ɮ+�SRʀ!?0xPrW��M@v�+|�P1��S�~�؋������%��_�����=&����-���n[T��-_�o.`��Kd����Z3�2�
���T8*O�ZhCSh{{֗sð��jf�ʜc�A޵�]�%#!PhG��'5� H�B٫�J�C�p������s��*��-Z*�J��h�����i|��L���yѽ+^�Ӏ�A~Y���Z�F.T0Q��'��JV�y�G��&�0��F�ş�b<6�X�c6?���i�A�ز��� �q��ty�Uc#FdZy	Jr����Ւ����{-��F#����-!LdUX�o'˿�1�w
��
4OM��.�F�7RP�lZ�k�F���:EIx���[�)�ۤ_��_E�6W&	�݉5reOD�O�U� S6_Ԛ�<+��$ �c"�M�T;��,�Ϯ ̢y3�?�Bf�0��di�ށKv���
����~�n���C{�@!�S�����[[u�?��N&�� �.��Q7����n�Ws�V��3��2y����m��~�h pz11���ݏ�}&O�Hx�B�P����t��w�%߲�-��~�䇜8�cOE��;xg��
����M�K-��#s-��ck��z@&,����0�����D Jk��U����Z�ns��M�V��Lh(������,Mr�P������y#�=���p4�z�ϟ���	�fX[R��������C=�:���(�Q&o����ZB��b(����<%ͯ�b�U�0e�R}�}	���i�b����d#��c��d��ĒH�.
��
�����dv{���H䷤`8j=I�D��f����h�cy����Q	��i���ӌ���}Dc10����l��]Dl�hW]�s�a�g��,��w�@�N� O�䥩��j����)��-w��,��.TG��6�o�a�����$�7[L%��q�S�Xd���YF.*�]ѩ��PE�[zv�_pp2��83i�3��/.]��p��P��O5ϟ�f�il��c5ʟ�NY.*G�raʴB�c��ϟx�*d͓�
�Ȱ4�w)j4{��q��������e�����4x�W�&�i�a7s�ʆ]ʲ� �ع��̘+�:G��x�x������~�Hv'5����)�v�һ����Ţ�%N{���C�]��E C��� �5�:�u��@���]�[4����l�$e��az��f�"����\� ttc�&5Qw�ߝ1��0�Y�k���3�^X<&`�[�9=a4�N�p������h��-�(O�����Wϖ���\TW+��tQD����XͿ�8���( / ����n���K����:/��H������tl�m��!��� �A����1�=�c�L��T��̵�˘�R�s�:�����A�,<(��<0�h�!�l���ᗃ[�c����18�Km�uq�P�
�|�g$�ua^`�n�9������)�^Y�����,�cy��3�$��i����b�#�՘#��\8��2P�Rb��QĿ���	�� o@[�p��V��<8
S��')Jxȣ�%��FZk7��W��(�cꇜ׏Ӊ#�IV+��;;��#9�J2O/��j_TJ��nbӾuB;�Bx�<��"<�Yj^C�EE��zU�߿G��5���Z��h�1�h�R��4��3[X�o2H�/%�o�����sY<C�i�����R���ыʩ�
1N5ꀡ]S��"P�Ҧ���nt���
�R[�7� ����l�+�7x�8*j$��6�U��2;��� 
_ג�Kj��(T���������,�ښ�|�?�n+���MU�}��i1���L>@��*�$�Ev	��B_��N��e-�41�����P�C(����Ë�ю�TuU#�pŮ|�"��0�r��}3,AWہ��&1��z|Y�ā��w�`��mJz%���	W��g!n�x� 7M���nw����XЙ�]Ҙ��o;��n�#�k�-��kT������y�묾�,c~~S��ņ\ݳy^>�è�d��G��U�+�B��CC�Y��z,�Ϲ�ͥgьyӧ+�}D#t��S����H�'n�-�ʫ���g����]>r��j�AO3I�Ǝ,���k�|�&ǳ�[)"wr@�!��^��Iu�8�2.j�ߠ� N>�x������ɛ�f��^潜6���:z3�]2�ܛ��x^����g���<y0��:d m���|��Q��v�Yimip� �u3oN�����(XC�-���0��@���Ҹ,���E�T��7[��o��#D���J*��x]-����Ѱ��؁;�����;lKM+��i��C�w���}|X��|��	��"3~�0��]g�bk�'�_Q�t��r�e�@%Q>+-�4O��������|�(�Z�J_o�RZ防�.o8^�O��r���*<�2��{ZS����i���s2�۠���ʠw��P��^=��1�_�����G�>�����]^�o����#�7���e��O?�T`����	R�k�жi�p�g�� �����Gt:˽)v�a �)N�(�0�w���]X�.b�taV�}	W$&�ܖ&�:�;�[z��]&]v�'�X7������%�QU��}D}Jd�Zv�O�Ν��$55x�eͩ�V��M�\�.w��X��
�L��(���&6����F�s����QW�Mn&���V"]
��������a���Ҁ�q��H�"5?)��?�rs�;�Y4M������3œ�Dx�,��y��X`�6%s7պ�P<aP��vю ��K���ɛ���,��3�����ͳo�� �����'��`�y�,Jc�Q������oܔ�o��H�3�����[ĤbC�=ls���G�X\s�;K��w
ǫ��Y��Z�gt��Ru�&���c�.�^�2�!t����s�nڷ&W8hF��!k�D�{�T �A9�Wŵs0���A�+ Љ�����eb��٢q��m�����iy{ǳWM���CA��΂x��ͼ��������
튿h�:vF�D�Qmʆ⒒uJć97/6q<D�|U$a�'BG�1iB{Ը�|gw2��v�ܞ(��TA�f���q9�����s�/ ��諺�O�ׅ��YO��3SƊ������~D���S���0h涇����z���M?�'�~g�E��YI��0Λ�w���N�Lt�^_�ľ�C"�W �-O�fǯ�u�%*E|��2UC#�U(6�zT[�4�G?�+cنz�u��h�(�!LX���s8�����(S������l*މ1���5O��^�7��2��>�$d��G;�������e��o1=P2�ZF^�%�&1(�%�'P�*��]��d�>BW�W%��#$ �z���K��$$Z��uL�T��l�Ȝ�/�Ѫ�
h���Žݩ$ �ӷ,r�zݟ�����3�m��4��yq�"`؀J/�n�mA0�#�8���M��PG�ԑ�\_���=�������BJ�����9�:*�ځ,���&Jˑ�N�1�]��ܫ4R����ДV�Ԁ�e񣉾��\&��$����Wn(��-����B�%UO��6�\#�D��糧�\�����C������P�)~ۗ�� ��|P���u�mc�T�G!��s��fKD:�f�8�۪��ѿ�d�<{=��L��b�>�;!�J�D\��^�iEk�R�������K8��6���
)�J������x�8#�P�d� {bhN	C��i��.��G���ƚ
�h�L�&�P�m}�Мd�k�ԵFv�)�ba��n=yO�`�V\�ğ^2�_/�W�1c�?�S0��iAzx��e���K��S*vŇ0��pZL� A�d��Ek@i�m�)FZ��R/��(Ƶvk��힏m��`�c�ܞ0\3��i�Y�$���Y5u���$uu��Wo����@��[a��G������!j}�s �S��n�н�|s�������vq�CD�v_���3F���J��f@"$���G7�e%
0~�d��!Sk��oe���1g�"��5g9��I�6���4A	���l��FB� �N�oLQ�P�e�`�1�JC�nӔ���`l"<R=OyiDvȣ�(�l���)
��>W��e��t�Y2���Q��.!�ڌ`�j�� ��������9�F�QJ�X�ѝ�P�h{hx5������/p�p`X�A\�&�'�Y�|%	��V��N�x�z�Eɴ!1�מ��4��X�X�}	/��&���D	����Ұ����nCE�K؅���X��ǵ� 9:YQ�M;�^���P{�04�n1�5����Eń>˨�2\��_S�H��(x��]�o��K.�脺��rk!���2�#~���:_��ȹ��c�֞/�^�X�l�����m}|�S�1�w�/�������uC!��n��\���w��� �`,a�> i ���`:��_��7C�_����#t�z-���Qm�i���EY+�Yp�����U9��--�"� �^��^m,���x� ��c`"�af�y���Xz�N�]N����n�4�if�L��W#��֠��5�z�ƽ�Y��F�+a��oܙ�8��;�G&�U2�
��c���\yj�}�X�q~Hk7E�o�h�� �m��g~��&);�JI����ދg&�L��҈��3xs���ӕa�̥9L鸳|v�+�B����7[�9�� ��"u3>}���.@Wc�=��Ʊ������|'Uk�5Aγ�#�7@��8[�|��8	W�S�H$��ݸ'�#j_���%���?G\�+�&��s�<�M�,�������\�HlEH2���xl�D�4]�i�t��	瞓E�	�MĐ�#�p@� �I�}�Ni%���F�B u@�Hx��T�{�N������cP���~�ҢtB��v2���v�[��iC(80]샵?S���`����-�ԅ��s��(Y���]kg��ԏщ\�����y��5y6�b�<'�_�Eq���p�sI�]A.0˓��y�j�fz>q7�g}��oZ�$�4��jʸv�7�:(ׯN�������{[� �:*�i��Ŭ�j�l	�ػ&��SƝ(��(y{z'� ���a ��1(��jC̓xN����pQ��Wƕ��l~= C�D䶏e"�����y,���	N~ft��C�X{T�(��=�(-(�������UB�����z"u��Bc����9��.s��:�����s��xt���Й�Z��~�� \��FU!8���ߢ�;��?���SW^A���Q�'O��P�p�A$t�4Z\k[&8d�