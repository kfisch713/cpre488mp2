XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Zګ,d���&�A�]z64�����_MG�Z���W@f��ا�> Qd��0w�E4�9�~ｲ*?�]kW�(H��'��D%&��_P~���J�OH�����|�T�54����_�3��!	X�.%�7�k)��V=�+�iVbH� 7]��rn2C�ާέ�����}�J�|� ����s����@5���E o��L�$���&��O�;���`���r�V3�
�L���L���H�0f�TI`��ΐω*����|��W�+�Fʤ%p�c'C�7�ƫ��L�7y{�I�u4OYi���^�A&��wJo� E��chC׷�W2M�Zk�64z�Q��:X ���F���v���I�ܹ�*��+�
�����4ȶ��}�c��/VZ(֬��[���U��u{+`�����^���䋥'�ֲ"m@�d��F`_m.����f�	]����X	�*{(9��H������f�G-(���t3�f�l��}ڌEb�#uE��Y�ȟ���#]�`9���cͫ��ƹ?�-,%���Xn�K:�
`�lK��/_�T���幊��헷��.y)��{YӲ]%�K�!�<9e�ڙ�ʫs�ј�J�����c�
y����־q;M���'4�svtW��B�_*�'ͫ�.���a�/��0w�&��~��Sx
��,R�jt[F4to�θ�(Ú�|E�Xt��	������j���"��:<6�yR���,	�C����<e��99�e��v����,�C�K#�k�XlxVHYEB    3d43    1030)�<_�9oi�V���G�*W)����q֫���D��na�CJ�$�.��:�E�ϙEw�� Lz�xfſ�sV��G���9�FRJ��@��~t�iu󣞋bV@���D�ű젹-
�\� ��Ԛ�o�tQ�?��1�g§�rp2]��T���1��Md���O&�|ܣ.��r�ԚR��L��U�G��u���U�#|Q��u�TÎmB�xibf,=@hRU��)�؊�c��JAP��l}H�r�2.s%�c+n�K�_��[;$i�H����Ԟ'�X�ga��J�8����nGA�]&�lg��v�8�R�t}�%$[����Ⱥ��ӟ>
l_�qH��3���\CQ�9j�&�_��<F;QY��������<��0�U��SAI��w�x5Kfy5��B[���wx��z#fRf^�a�"���g<��|�f3E�x�Dy[����?���FRF�ʠ�c���/y7�5��\bf)�p~q�o����K�]�t@H����@���(�ҙ��Yɨ�.�՞��'v.����	/c��E����P"��y��I�hw�c�mY��<�iPs�p��qz��{fj��_���@�h�;(Vyh,_��c�T�[�T?����M���� �m�v�u�M�V������zmx�pȢB5� �u��;��?XJ���%d��ZN����F\T
Y�<�r����z�����+�=x���Y����y[�����0Se)*��`�s�0��
0��iHbEѭ=ES��T�h�A�K����T��s��U���}߰Y~_Ǎ��+���?� ���E,����f���W��8��H�ήjռ�o3��p��>���kh�������Z��\�X����vIze��[]=��S ��j$;Ӕ̩<M	�F�QB����)��D��y�0�|��a�k�Ywf=_�f �lZd�����;��e�H�%�������C�%)�,�!	5BW|����v�h��$ G/�P�WV.\�B_��o6�^kU\?��9��vM�����2�ՠ%Wά�A,�8�'ᜨ������wa(�T������r6�V�A+d��8P[�rcZB���,�]�) �8�aF-��!ӿ�h�(mzU�1G���\��	
�Agd��̚Z1�P3����L��1�q��9���MԺ${�H)����*�(����/�>Stc,���iU)�}.�{�{�7�D�R݅�%-�)8����J�J2+`H������� l]=N��K<fV��u��\Л�nG�'�!E>�t'�|4��j7q*[q]i#�u�e����f�C-ڊ���e7��[�`���VA.j0Ѥ��m'�b)w��&��6E^(W�Ȑ=9�'�������4�{HQ�@�h�[�g��"�Of7��7(C�qD���� *�3o$C���V9RG���)&Wq��|ǘF��nvȰ�Iܺ�1���KQ�8��'H�:k����
��<�I����s9����=����2c���|��,�PQ@�Y���q6�-�,���̦��U����$�.��((�^N��u�A$ C�4&�z1�}�	D�l�ay"���=ab͋�~kmC�79%O�2POQ�6�/(=kLEǐ������*��H��\��΋ߎ�L�������i�GJ#6!~h��}�%u��Ct��l� �����p�L�*�z�T�ݱ�3a��m�1��������|[�q�y
�����{���	��t���%��-e�����Q[�l&-
[�<�e�����mX��.�y��Fi���c���r����K�%Fȶ���wy(�F
H:�b\�U���iM^����yFC|���<�`��_�ܥ�Q����Ī#1�����_}�~LPVb�9k,�ߗ:J�rt� ����`�L'���d���"��M�8+M<��_[��8AK�� ��i��M:���EK�N�q�[?x������bO�|ͱ�!�*Ȇ�N_�.�:��M]��b4�Z�cU��i���SԚ�i�
���fR���e���dnU����~?�֪�%E���'�;�8rl-xw�c
���i�[��- u��p�F	jά?�/j<�k v�g��rL����W�LS� �QrQn�`)u �hc��1KZ1��|�A�����d����z��8�����<���TF�
!��IP���JǴ5��A��ҥr�>('�ؠH�L��,�M]��Ap�3M_ 7H�n���,n�S�_�u��l&��I�*�>O����W��Z��ԧu�޶�
�.�A��L�#�<�5V߻Q��_���Gw�%֙���C�;��H�C[��^[3Q��j&��Ǜ�� ��ڣ�^ 4�Ҥ�ӊ�vb�n��r�f��~ �y�-�"��7J����#����x�������[��a}��W�eb3��`ȷ�8�J32<�"��J���{X���-�MV��;�l��B�ˀ�>�^]�ؤ1L���yѓ�[N���C�\fdfЇx����;C-�G$��#��;��}��[�J��@)������L�"TQI'��3	M�.+=�4`���H����������M��P#�h�uB��\T�;[\��VZ{v��6�E��5��~Ur�-�U��.��%ӆ��'�0�F����B�����85�Q�΁��L����[��3�g�ivX�~}^��e�����G:�WY �(ެ�,�d���wc�e��)U�8���v�L�m����]5cR~G�R~���h�zs�O߃��O���dȽ���}���ȥ牄�}#%2o�u���i��ߚXgy�� �A�WN� I��>���kR�=���zc����ɣ���J+�(eߥ3��
�M��M��5���*%��Л��mf�}�IF���H�K�h��4_s٪�����lT�������߉���G��^��`���1��*@ ��ХQ�3�	�c�/H�*ꩻ��ܬV��F$�v�=��:��c��V"f���`&#����9�{ـ�Uث]5�����6pb��tO#�Y =Ć�Z�n��H�����}u.S�
`�R�!���jԗs:�ޘ�L�M�.����,G���d�fw!���u
-|Ƃ�F�96�AaP��)X{��`��K^H$4�22��e·���}B,J]��c�"!_,�[
P�(c�Xƒ.T���	�5{|�_�����h�
"��X����v�F�H�f�U�\�8�=���d������i,�k���L�G�>G�Ƭ�z���U�2ѮlQ���:\Z)��B��A����X6�x���W򜙧3�gP��e�_z�D ԗ4�݉G��p��yګ7�4�k���x}` _�ͨ خ�Vh%��&1���{N;����n�8D,Nb!�w��n�����Q8hg�c�3ARg�D��'r��&�����n�#^@=�iQ�N�CCo�� ����L�7D��chTbύ��	��Cz?�G��	m>����ܑ�z ~UH�h�eC�>r훙�ck��7lddm�.��I~�3��?��0�28~6̸E�"D^�K#�����_i����п�H����
�ɺ>,�u�������Wo�ChgP7�J	/��M��gߣs�d��X#��Կ�v	)]Dq���Ѵ~lw6m�a�c)��b,rD+�7�\�_�c�=(�V�@��z䚎�tp����O.`����� <�0,A�}}{ق�\�~�ga��q�t����G��p.���P��@%��	9E��H��)�,�����j����4�܇I© ��p�\�XK���d7�0��Ӽ2IUYS�ka�Yc=47Q}��} ޚi��i��g�����M�ͺ3�r ��,~��|��3�M�qMA�̬�k��5Õ'��T$�3�,�9���������.�,$4V��B��Eh�6�^ q�<�B���;`E�כp��X�!�7�3b{Tj�������R����2��1�.���B^w8h($�/zSe��S���t&<h�Q�{x"b ��+*je<��g������{ڧ��+�]�i�Z'��_r��s�*]�*�)rV��O��