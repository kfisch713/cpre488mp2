XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:��z�[�0(��j~W��R���{#u���y^�̞�7����+��zo�Q�9Eݱ���;��A�Ҹ�Z4&M���o��r�\ �t��)�Y�my��'&�H1��L�F�rO�,�Jb�.9p����&�f���7��Z	9dͳ�_Gu��rc���E�>U�f���<LW��މ�P_I[b���l��f���#�XU;-�9T��䇁�L��(�uql�����&5*B�>��S�����%�h�ʰ�e��x�Ǎ'��hn��1ϓb,��Ɯs���zi�3�8x����.����J�:ˋq�
J�v�ؼ�E6As�@7;|�@N����r��8���|����g�o��p�Y���n�iP����h�Ύ����Ҁ��?X��`��Ӆ��J���&ʬ͖������1�qZ.'NVթ��3F2�A�o�{ 8�y�;�� �ri�N�h8�AE��>��E�2���G�@�V��d��p$~�'�����T
�]9��Z���͉~�_�ܕ%<^�yBp١��|Mx���c H��vr�l���,0b���;�l� �r:�=�g���J��q�0ᗣ��6��b�q䄃�˅��Re� ��L�(z��~M��ܛ��e�J��ޚ���/	�OLl	j=�wk��C����ͿqHzyN!ו�7y)��9��S��s)F�q�Gθ�����<��ߕ@r�%z�ǿ��TW����r|��e+e�wykD�t�r�-r�Hx����XlxVHYEB    dd8f    2160��7񄶥R/E/�����Ύ�N�o�,��N����:X[�D3�N�y�B{.@�ߧ2�����S�.=���Lߡ�J��.V۞=�c��S�����պ;��J���O�37���n���sB�����, A�E�G��\�� -��@�%�%�ƛ��4�����'[�V�h6�W���j���TwZ^�JS�M>���Tk��@��r؀3=��ǍT<;D�gx���q�(�?��QPB�?I�@'���^	�Uv�K�ԋ�3��B�e�3I0��4�=��k��D�e�#LI��lKlTƼ6�@O{�$��LNr�V���b������h��4�(#�8��t։ر(�'*�����z�{�f�I^5TT����������nl�7�;C&yl.G��I9ӛqч~���MP(�P'�b-�0*�Wqb&6gT��O�����_��y���n'�B���2{���j��f1���~��jx��(
�r:���l�B2�l��|:�᤟l��,y�)�'����d�l&%�ldז� Us�-��"\�G�ɶU�nkajP|h�Pm�9���[�ͩ�A�z�jQAJ#���bɅ�i81<�5���(���*搖OF'Ν����D��h�}��f�o��{�4�Q>���T�;�j:�N-�������O������Qj{�G�b�<��E����w�`�e�:*��ӷ�sh�ր��>%B��m�ZQ�A��j߷���z�v%�<6���7z��L����-�r�����;�2T|�?-��FO|kŲ20w$l�c��܂����Y�{ON������χ���m�� �<�@idn��2�ň"�.���Uk�~H)fLI����i�ߔe��5�W�L�nk�G�R��cǒ؄%��[<�}�W�:�T)��,�����/;r!D��ͳ�C�ǭ�
�F ��3�r��K�����ⲵ��\"��aw&�;3?5�߱�tG�N�-�v��B�.Qt�6x���t0�&�z���c��NS	Q���
��D;.:�4	�>%����F�7�KtC���b���2G,��mƼ��c;�(׷g��'ס�a���a�-�uM�ϣ�>'XZ�So,��ᶚ�����bwq�wb�����J$�wT�`���v_�?!��ySTF�
iˡ�؟�cϞ�dR?��B̒M�뒎xQ���S����-gO�-���ר;�����F��؀��j���m����lE��i	�1ew��t<)0K�#���x1��9@���w���g��M����N�ݹVlF�gY��	��:�ڰ� L-$Y�<��W�n��Qdq��E��0o�17�M����Lf�B��U�F�����ph8���ޡ�2h�%}7RC����l�]�	�e�W���">�N�.9�
�X��0�����H�,���c
��'u�޶;�_�e{$�t(f��)��is	�����d�j��g٩�G�C>�V��#1D眅�:���~^�s�kx���̛��;����v��\�|�C�Rx~��� &�#7r}Ѹ$r3+���Ŀ{w���~��� 䈻��v]�]�}o������M\V�S(V�P�q$P�/�$��0	��H 8K�p��aJXI�O�$�$����]��;�e�N�ԅ��.�h���[�<���)XR�`�c���ɛSB�7�~����u[�-׫ை@a�p�������'���6W��2� v94睊�R�V(B�7�"�撌����u��]9��'�N&U�Ɔ��E�Q�� �\���蒣�`�P�k#]�c2�Ѻ��WM�P�/F�n���!o��DgO�J&��$�ʮ�����r�Ix[n�/�|*P�F2K�N���β#���co�N�g�B5���wp��s@f�X|ZB�Z2�Ҁ��N��r���2��)0|Y����Z ��J2�һ<w3�S�ו�o5�~���h���{2��r�<i��~	�G��ip�\%�Ą��ܿ=:���o�KJ�3B�Li�GQ��hޠB����h

�����Bw����8ܨ�������>r���?�Ê�}�V|�C��Ih -�v_6Y�R;��)bx�v���x�g-��[�^��9�� ��"q�71/I�2��Ԋ��&v��&ͭ0�0B���hLl�f)Yj�W�� ��I|�;	W�r"�q���Ȥ�
	�8��޲�!g/��ԋ��;�ʮ��ndF[����YL�yS��x+#����s�YF������f(w\E�U�S���
�	Q��`���k����/�	��mR;3�e��sx�I�K�+�ft�wn���&�AKɋ#�ެ�����)k	�J^��2��]r�$+ڞ����iZ�h�Ğ�v��U��;)n�k��Q�&��g��	>I����b�b���#�A�t����ȲQ��W
{RrK旿�H���x��`��?\���o7�ћUz4�F$3D7��r��7�������}v�kSu�m�CW��Aw�}Z�|�-j��!1=�yMkC�߂�?��{1r�
J��.~I�C.h|o���1��ҩK����*�r$$�HBRp	�*��%+X[�.�Rl�{�����uV�o,:%��n��xTSy�ro����&���A��v����ck4� D���n2�Mv���@�ej.�`N��(ީ�t����WNLʧw$']!B>��g�>[����E+U�"%nd�h��+�0�L*���1}�N�Q�m������hP��i2�Y/t�o�*��Q=v��7��a,C�00�H݌��4�9�+=�X�#��)�*S/0���1�J���T�YS"�~�<Y��|lv3�s�Jy[S|PA�3v�������ȷ'�w��M���pkyp�(�9��t~��x�  vs�$��:d��[��$���E��aB����Ԭ�(���
�v�@��A�Q��Y)@��uXIcc\��4��F�;qy���?�*��W�ʦ��u�A�a1w���x"�}]��9��:i����;�����!�x��h��ǰ�^�d�R�*�/����/qi�������߷aifQ��K�p[��-�!�K"�_�`uT[����r�1)q���&HM���T��<�wU/��|��9����R��c���R�X��,f�v�.r1]�'k��R8��>�:�OM���X��`R&lH���&����5p��1g�L�Pfj�F�0����=�>8��9n�/�GY�If�庒v�#j�gA-I`}@Ll只�MX�!_��/yܠ����Hk�@��I1ٖ:΄Q?��Nk�<4oK��z+%͗���XY�5�����>E�����ǜR�ӹ]q�N�EEr2�H%:�3����n�g�n��)`��\a?�XAZ�5��ql*���#G|6v����!+)Jx�-���z�c͠S8��U���6� X�|p���D��54.l/� {Տ�t�tcx�1��^�`��Gh��7?�1�D�]��3	��| �U��I<;��0=��3�8�,ی�@�!O��C@�F�\��
�p9�L<���Ȁ�z\���|�!��c��Y]��T�hfB�?8�>:�ޘ�/�n#������i���k�"D�'��p�XU�)��������ђ�����)����'+-��}V�v.�&q�����1@�U��Op ��DֈzN�ߚ���`�8�gԓ��h�y����
��yy+� ^��DJk�y�Ξa"l���>�.$���8�I�6��eb��yI0 �s�Ԇ�~f������z(!)��֪[��P:M��f*J'@fA�v8�I0>��_k�>{��H�}I��lt���QK;$%ig��m4��z
�q��$�}�[~*VK��bQ|��.���7ē�B�@�<�%,�~�
��kލE�Q)SJkLk���2�J�J���Н]�3g��mp*�Ƚ�"ҽ�ه��"���{\�A��	��u!፠6���~0/�L*�Q�O��\_������(���=�g@	Y�>�	V���S���̜�U/N�m�*�w�t�]<�q�+ѝ�ݲD��j��]ap��~e\��7/�V��_��*?�ݮy���-�Ɓ3|�������c? ��,��>�N��4�C� h���?�v-�~�zq� �-�e#�6��C�I�WZ�5t�]���ƴ+nwa�m��,l��A��r�'�jޱ�A�	��ހ@�,/3���摹7���^��2ӧ�h�ź��L u50�+_ߤ���J���#����P��{r@�/x�Ƿ1��`v4�Ft21{t0�-RL�g�l�؆8m�?R����q���J��b�8T�l�wE���7�gM�V�Ww�W��j���!J�?��|�%���P��Ox��O�8wO3.����&�:� ��"4��0Qpm���?3p	"'�FO :DdR=�5�t n�Z����e+,Z,m�)?q?`�$��w���N�A��8e$<�%03�#G�0c\���\�>y�,{*��Nؘ䗽Ўp?�ۈ��<^~H���lM�OL�G�+ͣb�CM�g�UZ�+m�Y�����C7���H�i&�>/����a7*]%�4�Pu��~�5F���P�	�i���פ��[�M�L!�o�F�Ei�^	�N�[V�5�:��,ɰ�qZ{�m�9�A�ؙw�cl���x��X$7��Q�1�6�2*ȝ�C��%8��`#m{�`��B�l80�dc�攭�,�=9���Bb�'M�J�����<��-d8&�ڡ?ӄ�" ��!6��MC�D��;]
AnH�%��fd�=g�nHs�M��w[T#����Gk��y�	Ȑ_����'g�]H���~�e��!�Ja�F^Hv���+�0<��3:n���^�d�?��{dd���!�J���$X��|�Rt�'d��i��FJ�#:IйZ��~�W���8P=V����ݏ����[�uW,����E
�ǂz؅;��]y,�b4(�y�x	�թ��2 M��1�����4�A�}��'ܱ���qp��p��e��Ϝ���E�N3]�L=�yȬÞY�~_��L�!�xWI:a��V6M���WՓ2����<f�e�E����"�����Q|=5g��fo�����Vv3���t7��s�p�іl�h��d��l��s[��|
Qn*�a���Byfk�<��~
�IQ�}��J��o_���˭���u��}�Y�Yhbw+�W�����2������~8��c��O� 9��-r[�w��wN>�OB8d��s�3�?x��CyP�,Q-��Xf��<��ƒuY�$�$*TsI	�E�_�ʶ��Y�2�&�?^����Ҹ�]�oA��H��,f1�p���%�����<B*�#jǫ)Sr�ڐ��D��b>���Ч�{�?�8%C��J�d͆��e꠿>�LϷ��
��γq2�?���}����䰩	�Үv���'����Z �J�3#�a \6̵(t���m7Wm�ɱ6��$�����<�ʜ�Ś�anh�s����������B�~/�Kz��1�Iu�����wD�<}��G,7��m-�y	˫��&�;8�a�RL��r�и8��ZC���JtJB�[t,VۻW�)�gCw��rطZ��{���m��d�@ �H��I������&�ѫCS���{��G��ƽ|�EĥW�ra��0���7��{c���%-�i�&U�0��/m<|!�u��2�xWx@UV:%^c��vfV�%�1�pv��!I���|;�غ7A�D;�3��(���`����⏅���WO��_V�{��#wR��'ɒW�5�<�1�p��ҹ&����P�,y;�{���� ��G��Y@��E<~K�P<���g�v"�A�t{�m�~FK�ӸB:�vR���_]��L=�sy��֍iq:�R�K����͖��+���Jᡬ�:�$��yUQ���s��U�����`c������֜[0�)�}AQ>'��]ɚ��TES�$����ؒ!�)�q�ђ�o�t�{��Zo���Ui�G�?x/��ٻ�tLǨ|*���M��8%�k��a��=��l���P�'��v��W#J�5��p��D��t}#��UA���EtDݘ���U|v�(զQ1P�U�LE�͈�tTM���S$��v�ܯ�H1�K?
�i���+ɖm�EK ����$�:8���dw*��:TA��U�Rp�T�{�%�(����
VWs�Ͼ9��-�v�A.��f²wD�y+�ZG�y ��N�,�R�H�ooHH�M�f���͹}�_,��O�����LT��ဉOں�m���0�-��R$���=7�\��w�$�<��%A�M�9�Cih�BD8��J��1����;`�6�籆Y�(�r���зc��Y��.a�N�0��2PQ�o��M���~I�p�76`��U�~G�HNmE�TїFj��y��mf�dC7y�h����GJ�EG�ą[�Pcv\6�9�B������ơp����z+�@�~�����(����З�!wӌ쥀�ȗ�8�E�zF�r/��D|㟷P_PVd�79J�\9�N.#0��:l:�Y������L��S(KݪvZR�1b$ M���?;����۟��<��|B}�,U�U,-�f�=��!�΂�<иd�Z�O�ns����a33X��B=��g��f.f,y��ޒ��L�D��OPu���,��k�is9^�=�lW�l�
�� �_d�yڜ9�S��XWP��T�#�mf+�iҔ�ލc��tMw}t���3Ŷ�5�!{3�%�G�\�$t �љ�������h�oM�Q��|��}�f�d�5}Ii�6L��p�M^R�s�;?��(���4�[������¾�lp6]�ϬG����7v��A���Q�jQ�l�[��5h@���W��v�gbQ�^�<��ܩ�\�y��*jUc�]���3�h��0د익6*�^E�|DQ�x�V3�>���c� #�����
9_��7(D��@�_�nb	���;��i����F~����E]}f�H�MR��u��]�(i�,�t�65Zi������m�j����60�};G�?��v~T�-Ls)snlyg�'h�;},�7S��{v7�e�0�w�?���1#p5�>���|�W1\9,���� �晎Z1Љ9ac���6@�Ŵ%b���5W�i���wJ7|'�۹j�,�E���W5�"��r~H�:��*}1h���ae+V���.E�gt�8'+�Og��F]}U�Z��tw�&HD+��-���o��+Exd��156��5� ��f[��j��@��i?t�{�3���t��%�qNt�=�ڴ��U����~�&���S���ײxC���2��.7vf`X��]��/�3
�����Z�6�	������׶󿡳���|��Q�u�G�3�B=t�R
n"�GYL����k�����?Ƌ��h7T�{Ƈ$�+�i6�y�rÓY��8X.��ɷ�:�L�����0V�#����B-C��� �ף�'^�>Dq���*�!��&�g�6�攍�zqxb��?�!H$PHd�C��_�	��s�,���H����0����j�дdf�l/��M�_/�̫���\L�/�r�� �Z����� �cS�xƋi�pv��Ty�G�G�yG�,涭W/���V];�Z����4q����n�I�	��� ����<5D��u]6ҟ?�)�-d2�L��݃p����O��PW[@�͖e��zE|z���R&GI~U09�Z#oɫ6��Wta.�=�X	����vq;�>1(w������DO�B55��u����O��'��YP���-�Kn���]$����]�jXy'}�	��D�QЯ�E��^�R7b�ŗ���J[�x#�?��sb��\?x.'�M>k��.�[D� 0=�U"L愁EF+�>�X��f~���(�&����8����hU�U��.VV�_����2ܮAP�i��~u�d�����5��gċo����U���@3P�@�7�ҞyXWA�K����1��c	Y9�eb�7S��	A>�hz42S\��B��42��9�Uy�:�h+�rX7����X^k�#� C�V�k;�a�e�w���/+��}�����Xh�8(�[8Q�-6s�����~b^A�? �5jڅ�� ��fٯ�\<#����!��`'�84G�n]�X��'�2E(`L����LG�*=���8Z�s	8�`�I�I�.͵��Q�U��!\F���,K���a�#a�$�/�r��_�߮
��C�x־j[ƪ@���C��P[(��ӵP3�uE�%��`�W7`nĭ��CV��	�;ǉ*N�RT����e����
�2�� ��8k��í�kդvI��l1Wt�) E���l��2=Q��D�S%)��C#Ud���1a��^���M.�珗#$�Ay�ۘ�