XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���vv�AM����]��R��"�%��H�g� ��qS�d�[0�"D�+"Aoj$+�%BC�zG&�3�}	��"��q��<OČ��̼�R��
p�
��[-�7�pl��J��W��sFˬ�%2��k�?7�����"`��5$0�I��32���C>��U����'n�������RL�Ѹ|AG�c}����/X�o(��]<K~�޹(\Z�ʮ@�LjPh2�b�r�]��\�S�V�B���;aI"��f}'/;PC�|�KY��dQ�>����ZQX�.=�P5�ir�H��&������4(!la�E���&("|ڍ:�_���_i�h'����p��2@��+�G:��b} �ӧ�T�ȗ��5��!t�W���Sf/4���@�W���I��>��� ٺ���Gk�f6""7Mx�5��\���!�ּn���������?:�O�4�(2��P�����Nm0�_��k�����������+Z����k����::�Y�ʇsї���:*��!^����:.���B�"_����b�qV� �
i_�a	��A�������§�WQ*�x�Y�zV�&:O����������ev��6"[oqAܵ8^�a;�{�ꭘ,�s�(�J���e���ȑ[1���H�������Q�������V�&oW�dm�i��I�b|�W�BuaT�_m��D� .�4���Lol��9��ɯ�2�65�Bݮ��k��h��U{HR.��v����XlxVHYEB    1a2e     8b0&�@^�Ⱥ���[�s)�T�/H	vV���w�솗!�cli�Y݄�\���(q��I�]�3t�jn����#'R 4���f��rX,&�m��N�P�y��⽿"��n� ^ �Y�l|{S�@����%��9�56�_���횉���hN-����h�; ���S��15.�����K���-�<��c

�E�.Tntc��.�j��Ɨ	�&�s���OC2�	U]�%�͹����g�jlŚ�Nz�������u_44=hj�:��G?��r�~96Zg���E�>�c_���qEd�E ��c�K� O(q�]��&dS/QF靑iD*�wnuym5��J7BA*���k��b��'��u�����������ϥڇ/�k'G?���,�v�*;�a�~��FS�z"2?�f��~iݪ`�X8�����e�nxL�<A�S�������a���	P��G�4����F��S&�|���4��
�z
n�e6eo���"R�Õ*���6�3R7�ڟd����xB$�y�cq@�&������X�]ͬ�NO,>%^�f�gń�S���QC�Hs����T�߁�.��?Q����`����Rd�����j�c��b���~���d��/&��]-	"��v��@�3V�P�dm�o^���Ma�l��9nz0
7������Y��QOΙΫ��^��U8�~��#��5�Ѓ�H�I�;_��(;b��'��ρ���$�FCGL-gVw�n�ѷ��i��E{��)���w����)x-m�%���'xq��I����4����g]�SJ�4�؜A�Qp�I�y���N96Q���Ѵ�*R�s"��} p:
���h4�}�7i�%��rd�ƕ�5J8�Q�?n��ͧ��W�H�W��O�������c�Z�����E�}�L�s|�I���#��8hiL����zj�>需v@��k[«�6�+|�a(j��]�����~݊F�C�)}È�ո�k��4�`Y�y��=�T��PS^�%q:n�/hЀ�����@u1�VX#�\�aF�9�4A�3�K`��+� n����g�'�
���u+����7��jj���~P��g�)�`>8Q)��{��u:�W	nQ�A�ޓ��:�3�r�$��3+Oa����kL�G��4�qk���2SK/[<�=�	ݖ��`~�1F49���2�w������9_��Fe�}W�ts�I��gg%�N��*�g>�ާ��H"S.}��_��'y9�N�7ѓ���
�S��PzD�"h�"����;Ri���m6=��ɳ_�����#�ވG�0ވ����-+Ԥ+P����I �b �U��\w���JN
����l�X#yw�N�l������x�⫛`R��:�5��P�»�\�e@���8U��pޝ/�C��CI!�~�U���۱��-'�b��|�ƅ�b֦���lq|z:�h�{�6m��O�I��+�S�2:&T:l�Bl���`�C0�6����`�ٝ�ã�m�B�'� "Z5��E�Q�U0�ڬ��6�����g�C��bH���[��ڽsS+���W�Vn.�´�<� ���)V�;Lɵ��	�B�i&�P�o@��7:^�L%ǋş� ���	~_�R@�{f!]��Z��|�.M>P�b���ˤX�wV����>Q�:�n"�0y�6VO�?2݋�g�<:�𻄥�+vV�� w9w;EA(5(�j�?_��+&�Ly��Z~/���I�79x����p|&�9�l%f~I�k1�;Ia񤰉\��"�� ׍��JK��j���%߅�_�V�R�:�i�jE_�+L�9�'1��.�4�q����w�ㄿ�ƕ�XD3Zힳ�*ӓ�:[��@���tO?ߞM��o�b� 1G�_���	�	�).؊�T����7i���xۋ��R���=�CEWLV�G�E�p�$�K�z���MO�QD^o��z[���rr���ΪB�֋m��8�J��е��񇧷��ף�'� E�y6_F�%/3zaV�	R_'���~�u'�'u�sd/+��h�	@�
B�YR�mNw�Ep���j蛘K���ބ�ށFȫ � ��C�({,�G�8s�[u|2Q�o�ݭו�^�;
xN���J��c[��b[����HjPy�h���u�܈��PJ�P