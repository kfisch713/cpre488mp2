XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����E]��U�U����P��Ͱ/��a�<��Ir���?�(A��*�s3j���Mr�r�Ɖ�߳����CJ���2�8�����67��j����ϯ�-�4}<h�,i�?�/'�VL��16�U_5�~w�Hd�KGOZ&}��\�+��X�5�->Q��~�h�=��5�C#6qz��&��U����9�4��m6�%V;���D0f����Z6����8E�j�= �\g���v��c��UU)��b}ꝺ)x��o�,�I�fJU�9h=��nh?(�L:�h�<�NX���_���*��9�l��������S"/�'|�{H�h\ait=��Z3����Y��{Q�	���s?$׃J�͒��{]DJo;݅3;�K�t�E��M�p�{�հV�G3��-��`N��8�3A�����OϋX�Yj\0��XTF_��L4�G9@(����f��f	ě���L �� %�Ԭ��u��3�.���O�4���8ഠ��C(�WN�87T����q߸F��2��Z1�jr���b�g�s�ٓlVM%O4�Ŧw>	��l�v�t4�������R5��Ϯ�\wx�mmh��^�׆�z��'��fO)c`6a���j�������RW`�LW�dZ��7��U�¹[�9��->Ѿ�J��fn�M8�֤76�p}�������#U�ri)�4��6����q�qM�l��[ɂ�j��qŽ�	w�G���*�B����!��x�_?�p}'�ՊY�BbcwpY�XlxVHYEB    6315    1790Jd��}�%���#L%˵~t��x�^t���L�K$�;)��=�J��G�"4���U�4�G���#&Q���0/�38�q'����O�*"S��I�_��3z࠹��t�7�j��V�}����'������d�ȍ�zb�����927��{p=�9�D`���dm��1/�c�U:Y'0���O�Ӹ��I��� Y���M�9�*�yo<��߃8�?4Ѱ|~/RB��|��AJ� 5h�ms�����Al�������8xiA�L�c�5-�A۠����(������ށ�+3�F��L��ͫs� �m��_ʋ���5�j���nun�F:& �f���G?ݦ�A/3)��h�N�`&U�2�3��4q�1jXv2R_�;���}Y�'�}�6Am:7�'}�<(�\X�O[���9G����oMp�gWm�{���w�2M�����ɿ�\����b%:���y������+�`�Z�K~�	����p�C���-<����ʸ�i�h���%��_����2|Cs �z��D9��c�?�B�����_�-�bW7Y~��1���oֵ�+V=����ð��r�lM�]S�3g>�H��z,��-V���c t��O,[���I�_�,5��l�Ќ�|�Ch�m��d�4l����1��y�a�}ю� h�i|s0���/�%t�^F�梷�;y�f�0N�of����p`.ax���3,Ɓ�-�y�����U>3At8ft�'1���V^����#{6E<Y���u�;w����ó{
��C�[�c7�bM�4�S�_�>%<t:��*RS�8�͂oិT�~\6y�p�p��j8Ĥt5IDn�D��:h3��a>Ï9TƔw��v���H1`�E�ڊ�*ˇ=y��w��W��]Iu��u����We��>�s�[�PxJ͒ṡ�4���[!�|+�s�2Ց��Qf��IV��Z� ��ʅ��~=�->�.4D$*�JK����`.e񥶱�g#�����j2�E=�Ѫ�I�ȧ�#S'0+�����#Gc���[�p�f�[l�÷&oOP��,�&�}��w��8�[JDɈ1���>�ڸX�PE�>��	��w�>1����ϐ�r���>^U�'MPb+�.���_"�$�=�%A������Ȗ|$�R�Tf�Wȟ�I�G�mU���͌�͜��t^�z���;�l�Z3��(�8_a���q���|��qq�6�5oZe��5jAf%���)�IJA�&�ʾ#�PWk�g��Z����t8�*�`y����a~�&Cо��jz�ɁJ��
�S,�k(,���+�R]2��|O�Ux��'4E6����`e���:�Z�5	ǲ�K�cU��̲����|m��O����/H%�O�Ov��<by �}|a�O |�l8ۊ�M%'�,�V��z�������0m � %-��Cm��q��윱�.n�!i��>$j������ZAj�]��F� �uy����>/D��UVk��Z^wYX��EHR���"�|��A�*l����9ɬJ 7�F�1>��_f,,���_ ��Qi��T�d7�d���30x�V�I!�v�P;�Vo��z*�X5��П��b헩ʪ�w \��0|���Mn5��[�]�x�.��O�oX�X�p��Ћ��q�J0c��v=]Ź��3�Q��M����Nآ ��0��x~Wؖ"�����?�E7����4(.���q��Mc��b6�����Ze}��l1�����h�"�J���d��<X2�>@j,Ċ����Ç(��#�a~�}��
zښM����j7��#�<�~.T�0�v�p􀢁9S������Z�U��X���TӅ���%е��y�:�A�}"-�d��C݆�~�5�"x�-祭�l]���-sV!7�#
l����:	(�ڥ�F=0f�%�����k	�cj�E�����p��h⼞]q�/#~|>qqEfR>�>�	���	/`v��5xZy|��� dgX7��ԏ�|���_/��m����M#l��M�;�WPӷ�!�u�\A(��~	P�F������k�Qg�����r�Ϟ����ß��Z�|v��4X�-�><aO`fá�ٟ3��6���X�}�܇+�A`������]r!CEf�R�I�]�G
����"9Q���x�O�uP���mP�v��	WP�����Pٕ����E���T���Cv�n���u�9a�1���{�gz[�>u����x�%B敏[~���B�|����~9��Lh!g��������Q�{����JSF��sy/���k�5�4�&�;z`8<p�>|�&��Ì�[�TB�$؎�8��4%zo�*łuz�ާY*0��gRq�!]Y��/��f� ByLm\#�-QP�qN�����ܗ@��50�D�*q@J���`]2��I1*��s"Og?}	��z��y�(
�B�H;���j�\2Uլ�n��
�8���gcN(�m/+v���7�����L��?��9�<}��P��´� �����޴��6��1ޛ�dw&��B�]��qv�ŝ
%4{�ϊ�.�h+����Jn���ѷ��WL�ь�uَ�m�Lvk�\n�1��O�3�4���i^V����'`�rr��PX��^K	9�s�%H��Aɓ�T, T���2�Z�: �Qz�Ų�/.���d��h ���c\���P{I}j��p
� �$�;m5�����a�&�s6gU��»'�iV!vq�n*P5��2A3գp�3����h��B�u'�ϛ#�IC{ � A �jmD��*�{lqzw�}�#u��~�)������>b��S�r#O�9̇�$3ր_����l�mVQVC~��z�J��8F�3XgM�%n1v�xHFh(}ҟ��'^�\��v�+�"�E��sB��/�Ϳ(>e���AK���I�p6���xj8pN��I�岢{�:*����sŨ|^��y�ã�"��ݿR^M��H���:����*��e
b�0`�ϽҰ�lG֮j��#�"^ة�W˖2���YRs��� �Ǎ�d	Q��'�3�csL�`�\����a�),����F�zd=7�b'у������/-xO�8X9���o��8,@%8�°��>�8�'3��B
��1�ӭ�T�VݻY����D�nc�	�fb�"�\�
�, ,��j�d"������u��cK1�AC������w��8L���ޟ$���8�e�̿���h(�ڥ��KIE�Hf �7�o�����)80�_	.��/��Ɋ ��W�b�|S�b���D�����^���(�a&�f����i����@�W,ǂP�]Wc��J&b{h#�E ?hUC "H�ޓn%=I���n�!�
��5���E�-���E�+6!��D8,M��$�j�V���5��[�8���v��$���p�R$�y9��|�ݘp(V�ټ~9�3t���&�|;U��6�>��j�+��ġ
�<������.?�l�<-��g	�	6�j<�0���c4�7=���/�@R6�QЇfg�_q9�4����ng�Ȗ.�8GO�|d��:�o�#�hrSw�w��ve�wW�k�a�ߠ ���
��km�BϻƜ9G���lϒ�SV��	s�y�X(�ډ3+4yQ��o�|/�5)lT��/�WWٴ�<6��`x�w�e��1�uc�:�������{hK3��3�%8���?#�Vl`F��m<&O���"����� �d7�+-2�QB"�h�B%�?����5��I�PA�3�jKP1�4��Dq_j�O] ��x��1���Y��x�0؍Z��@�k`�<:!X⫠9'D�j��Y�k�6b}��[���E7Z�Up��I��������F�:�\ˇ^&����p/L�����w��Ӕ�Bݫ�Qv�)�.Ԓֿ�"o�Ȳ�fH_�
�Ug���h�=���9�?��5���'y!|S���~��飨�58�)������/;��c�S��L"�jJp`S��2�W�U��Z'�R�x�I
��3O)[��!(x|��6�-\$"Q�	ڞ��U�t����i���S`"v?�\���J��1DX�M����_�O���������Gpڕ˭V�K]��;�X3\��lvI���VBT*�L� ���'w���N=�+v7l��� ĵ'�D�� $�;)ڱ
��)#���?��5��~��#�y8z��
�9|��e�����P.hZѱ-fL�6ׯ.�?L��^Ya
W�N��l�I���j�wH�#JO�sKۆT�z�*�z�xpڷu�#�:��uga|YV9~��'�)X�q�	|!�Q'Ȃ��Wq5+�������SF��A5��s�uA$ܨl��Ѹyl����}g崶��#�'Y��Y�����E�ƽ.S�!^��р�_�I��W��\�=�|�����O�f�����G��_F	��Y\��^�|�]>��:^��i,�P�#R�%��nsEt���4��v:�������D�x��u�����t/��\f$�Mu�ιC�����A�m�I�틅NoJ'�>��rZ5�I����j�ѩ!�Ƨ�O��4���ƻޭ�RL\����M����B����y�g岂8���4�6xP(��[�9eI��.�o'hJ��[���M�G�b���gJ
^`ae�ل��ʱ#�vC�3�ie>�S$��`Y����v���z�&�t�c�8���#����]DKb)x�*�3����5v�F;�r�Q#!'�u��n�2�#X��q�cpx�"D�^����:*��J�˥U��f1U�w��F�� ��	�Ul}�X�چA��)���iؔcX����q��b-"�~E�P�Y��N*lI����'��S��u3�@�������=l�s+��X�U��1�u���H��v��H]�i^F=�B��x���vC� 󻂐#�214I��AP����� �L���T�h�C��u-�J�l������E����'��ًWz ��IW�6�* ���Q��P�I�5�_� ��Q9��������G'Y~E���ʆY�Sf�O�ᱰ�w�HAU��W(Ǵ�4 �fo��q�q^-^��]r��d�̬Z"܀�������`������.�*Z��t�#���u��+G���b��$���!x�\���D�GY�M����'��5��cH�u'��숩p/eb*'���Nyg��3Ư�p�r���<�[]�#�r����FP�ݽ~�2_v��+�2ƕo���o[��p
V1<#κ���zl����>�&�5���d��ϰ�<�����ʡӤ=��L>�ⷩ�v��p���#Z�!3�{�U03b��lӴ�Wr�Y啃���+%�N�pk���^wF��L w�A2K(r�DǪ�̘gw�r0w��@{&d� ,�iS��/�9X�� &)�>W!�`Ԇ(������x���fv�C1g���ju\}�d�{!χ͵P�?x�������\q"�|_�_i�
Ź�B��n���r��4G��m�r��� ���*x%{��4�{�Q���3+pdcE�T��J��dj�v*����<Κ�fl_�t�e�o�u������+M�p�I
���i���#I�#���)Ua������8���șQ�y�B�w���Z���ܬ5ѥ#�Ѳ?�����%ۿ��4�^�_��{%ړI���soڶ:/(����2zr�l�w&��@���a����U�3���SM�n�ry?��ö����>
��!�Q�7l�~�W.9R���x-`���I���g��`1��U*��� g��w>�T̠w�R�'��`�G"�r|��jd�@����k㠻�&Ǵ��椂��;�F��G��C�VD�'�E�,�������/Ƶ��_.�DV@�p�3�]X�@�a��T�� k�sȲ���'`Nk���g�,�h���?�`O#���.	�w