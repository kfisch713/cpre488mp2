XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[�0� 6J��2�{�ȟGѕ���s}p{d �(f��Ds��^ߔB�2��+��}e�=����` ^.�/':<qG��Y���~��n�Z�(~�2SV�Au�w�������V^̏�d�G���J�@|d�7Ax/���G�*m��¨������E+ڇk�K:���8a�b?�<�tƟ�n� K��Xt=�=��S�g�ꉆ$_��R~��,�LفwC��P6vs�����
�?����<27J̍>�RTt�R��5��z#��_�Y#p�����k}&�_�,�k�M�
Ã{�<ގ6��̖e�)])^�'�[��J��vca�	�߽���i�&)���ږR� r����E�DOWw���q��G�Jg@N7j��}�1	s$��؆�96�f~w��v�zȵ%�8� ��2B�i?X�=e�`X�=)&��3�B�(}����>�1 +F�"�Y�zJ^x�e��d�To�u����SI���Q:��>�l����\���[vJ�mHw;����u��$2UV��a�p��4�'�en��h�>�����ɲz!=�T��P��L�i3h46�c=��l
پ������L�6�(of�ѨV��a��&.{�oR��T�Xf��%Yrk�Z6D�i)<����p��b� �i������xޜ��b_.鉧��O㜅��Mu&�*:���ɥu������G��s��Y|�%ń=�UL�]\`[�vY�I�i3�l���}��������E��v�R�sjyf�Q�ަXlxVHYEB    95d3    18d0���zÑ�V9W������s㊹�<������r'��@�"^�a���t���(1�Q���i�3l3zeG��,	�b|:��v8V<�׋�rsJΠ�W���؃kf��O����ꄱ3#8Q
�Ϊ�P�9�d�� �5a3�>�@�X]�/�G^ſ��i�^d}���v�����B%���+jJ�&e"G��Y�{�2M�j}Y�Ջ['- �$�Qހ�r�嶂A��_-.CCtmG;���3R �wbvQ���1>�}�i�W�ZM���'�{�uj�J`Șv� ��e��C�QZ�\ �4�$j (:����>D:�9�7	�|�\�'7`��
8�5��}m��ދX�
l�#�@�N�g��I��>^;n�r�`o�8}��Нߋ�dK�ەvr30�J�������tiM<��ʕ���5����#��Ju�臐�@��r{� ��)ջf����n@')���3A��X8��u�6��>}H�ΣH���E�zÊ�	k�-`��]S��:zz����I˭�f,������T�� S����\(�@�xKFZ.�&R�=��F�y�S1��qN�r��_g�'ď���h�Pi/�/�ƍ5��;&C��ҽ��{����;k���mL8s�ޓ~#.L�yD�'�h����i-�W�ux�8�ϰfc�_�C�^�?�(i��F�q>Τ<m䅝�z�-)W<��B P��4'O�~�X��)Z�b�n|M�j�|럶�����h�kq�G���.��$�]>%�I~'����j#�>6n(�B�hl�Rp���$D���<��٤��9͖��z���Q]�F�OC�ɫ����E�����弄8P�q#$z@ȑ�3�{tP�?,���!߶�I��2ά��jk�o���&��F4�܀̥϶z����.���-D�^O�1�3����|�z]_��N���l>t���Ԟ�U���RW����X[]�rWj �K?����]]3^Ss=�}z��2�������S-оŇn�0^,��U�0�V���y��qz��gC�w��,J�-}����@��Z|i��N�Q{��P����1��vt{��P��.٬�X}gkÅ��V墣&h�ױ礫�P�i���[ݑs�!$U=	�P�<5��Q��H�Ƭ[k~�q�y'(9C��|b��&��ߐ�I�>L��r�\g�7IU�d�����~����7�c%�����"��.H�
 'XBJ�v�;Z�^�@��2�-�<����蓼��Yj`aĈ�RG��T���;�̯�*���	Y���j=
ROS}u���ڔ�͘�� V�Ϻ�W�(f��c\��aF�;=c�b]7`�Y��q�ī&�
 L�4U??<[`X��v�F�-�9�*�o?L<c�Ϫ����}=vc>�C�+�UY�\G�^�_�5	Z`�����e���M����L6���[�����,s9�2�üi��C�8-$#u�J���K��?sy���W�B�;w[ݑ����*}r[\<��ű�Ⱟ]VLiUIÒ�b����:7��{1
ș��H�S�m�Z�)��BfCǚ�	���hL���؃�/k}#
��,F'%�C����pl�)�?�$a�h��Wk���
e�=�df���
b�^n�X����fE٨KUNz�-���Q3r��NJ�i\��������狜9�X�m#jn�S�h��Ek�����~>��i}*ׂ	�>w�8��َ�R���I�i���єe���L3&�=uR/i%�{eY���sD��ҒR�[+��w/��F۞_]+�u:1��5F=�Q�A�����?��"U�*7�S�S9vF� �jT~�y.��˃u-��%�\�~��{���OU��-v�D�dWlo�<��K�O��_oe��w�Hc����Nf��9f�Yd�"��"�� ^�:���LQ�ҢA��fU�&�)��o���Ǯ���$��	����0���s2gB�כ�����z�ɯ�tЕ�{��aBp����je����i�?�{ݙK�/��T����5�Ķ���&BFA%)J��'���V��e��֛X5�#�k�ke!]w�>�L^�b��h������W��:�]��K��xߞ���*�)�GyBn�:X�?h:X Hh���܊�ط��p���Φ��Î�I8~&F/��4�C�+��`
��z��~�>њ��@��w�b8c0�Y֕�	
��&;��p[��Ǵt)��\��T�{8T��p�^{���h

�,��?�M b:��Q�l�W���"���;9�w��%�8��1����#��ymu2n|�N���-O�䵒}�m��#h��*
��I�*(J$k4WK
KβPrL�1kL�^=����5��ܸ�;��H����/��ؔ1COE�f�l�Q����3	�eB*�V;�5�J�>�FX��P�a��>�9 $O�3M�/�.��:\/N�_��)3�K���RaE�nX���QS��oV�D���B�����*x�3�h�mtM�w�
�>�!5n���/*�F4ɬ=�N���'}戀Z�?������5��Ǎ����ۏ�r?��Ó~x����-� WH���y(�ͽڏJ݄tMvoQΕVg��B�s[�Y���Sޒ2yjQ�Owd�Y�6��B�e�� �E��ⴻ���� R��?M�4h�ұ�Q#&:�j�����'���#�������~r���qPs�i��1����H��O��Eɯ\l��Γ�����tTn��v�x\�$?��P�a�VV%�����|����=��o��)E�/�������D8�#`[�Z����̛Y�z�g���\�XQ�|�� OA�����e�$�n��Wor�����/��<��Y}�B3�:���m��<��M����zfo.���4bM���e(��]0���(`���i��=���e�0�o��k�WO����Q�L�X/vJF�R��F��η���d$3�٭�U}��ɐ�5�EY�V��z�"������e�aʻ��zRKf�bmdX��9<����wA�8L��4r[�w��q��)z�ܸd�k��Q�[c�y|	Y� Sz��`�6���,�}���a ��FKm����&;geS��|�����W�5�k姲y���6����KQ+�( �q�}���\�v��E�B��V�Ω�O�~��CX���1RP��՞(N�o\�����	�����t��1l#�w�M�@��P�d�qw��y�G`���Mehy��3I�NxwG��52�(\4�_�)j$;ޟ1������|r����3eC�>w��,y2�ʜ�w��2dϔD&��)W�Q�J6	 ������'��'����Z���j���K��46
*w�~�ܿ	P畝��Ǉ�������!�4�ь�ŉae��x��_Q��^�4؄G�ɋ_���c�^.��I,b��w��r�X�h8�[����t�������68!�`x������2��V��/k��5e����x:*�7i�ͧn����P��
����g����&�����VH{Q�_��ϐ��#g�/���zz�q����wyF@|�����En� E����VQ�<����ƺ���-��n3�V�f��_z��q����
��U��Ē�����3So�!s�}���le�(�� ���lOw�ۤԼHʘb��B�J�dB�.YT�̗�Iڰ�p�6Vt�J�[��))U��~Uc\_j�E:�"J�xb�E����.�P�0��tc�Lg��2���"�QB\�D�o��w$*�����ګ]9R(qR��/�M�"@;�IJTzGI�{��}��.]�>�U��IV�7�Q�y��xl@���M��=�'�� �zO�+�g{bHv��ȼ��=��9��,09�ʤ�o@��Y� s~�&؎߽��HDw�Mjs�t��䗮�b���2T8�Rv�H�{��laH���`�8 O������T$����R����4�� ��@�&�M�^��[?����e�����͊�;$'-��I��jk����GL3�i�<N �pc�I�E䏳+��A)8��8I �@���S' Z�<l+
�|Qc?ř�½�G9��D��:΢�q���)�{El�$;�]ǤC���"_{���D��"�	U>dl�Ī�a܅z\#ТЁ��`�p��6�$�|���k�c$�щ�P1�j�	�����P[a@�bd���J�S���%M��l`��D2�(]o�'v�,c=d{&�$��sd�l_<���MW�*$�+��/�"ji���WKn�� ����t�)#��Q#2�0��z��� z��u+�g�{l:*ͭiL��7s�I��$}�W9V({M�عU��/�*uZ ē�k�C�@�(�~�I��%>êP\-p�W͹��u�}���>}q����B>�ٓy	�[s�*���2�Џۯ��l���1�Cf�˶!]M�a):���ɽe&v��/��h��epd��_�`Y�n��
��Gn`*�s��_ıR�������3r0��o��:n?�\� ��������i��K�\>�AZ���`����x�̓��Y�~J��Mu�����SR�È���(��F�t���VuM$���H��8C��2��=:�6������M�C&��I�,����
MǴ�R)��������ܽ_�~����"�]f(zq�oK8��g���ɹ[���Dwj���	�������\:c}��U�M-�t�P�b�����X^.)F�ѹ~���H� �T�-'ڏ�T����I	+θ[g��t'��\��E�W��VMǬ4~@�ɧ_���y���_ ��(�Q^�S4��@]����
b� 39a�`��4I�o��$+j����@�w����T����n�ӣH<���-z8ðB�ICR�6{B���	P]}�6)�����7�.�������v�{��}|c��������v]��ӏm=�,���r��Y��5�A��"�>sݳ4�̝�{���0�{%�i`��]���D���׾���4`���Ū~Q)���K^x�=����H�0L�����z���3�ge6"&trz�G3PcU�h�y����Y���!��`���9����'=�|2�]ڄ�>�k�2��ؓ�N�A����̏p3�����x�"��O��Ʊ�2:+\����#�-6����S�l���=gk�o`2�A���Ӷʮ��8�$��W-��U�ح��n%7H8�Pd	W��ީ��)��7�֠ #D`�%י���{��Q��2�ﰽ���U������D�d�a�7�d]-gZ��fpVy<��Q�3�f�+���>��.�hĐQ��!�-�}�_}@Iy�s�!�?�,.�Vuz��	0��v��H���Ս�0�{ˏ��W=�k�kaޘ�7n2@��͍�!����n9�J�:P:ϛ!N.�
��ϧր>�kZ�i,a{��V�F�P+�Y�]ԇa�R�I'�,�#��?9��8�֋�ZMj�	}�J���g:�<�\��Q!O�ZR�MSѷ����P����a��m��5����)�_/E����͞ˤt:=�+ˤ�κ�+�G���5�9���l�YN����&���X�H��O	�䴓?��ca�JK��nE.TŪ�C�%D�g׻�*)��U\���|���@ۥ�H��+_���s�=;ءM���mL0��͒7���O0y9˺����z��*�a��-�X��1�"�����d��S%w������O1r`�-��q�W���ۖ=�N�h�6DvV�'�8�'%1��򯇚�N�����[M.�F>;Q����t�|-�U����+������:a�jv�]5��&i��N���"=��/��^��:"��9b<]��Z>��/��L�k9��[S���?�[QF��5P��
�op�w��v��R%��Ȗh��D3�0��pTT���mK�aj���8��x�9�(!���w��F�].o."r^���Ǟ��{���[��!j���TCh�	B�F+��RXs����84����4�q�,��D�#1��������Fhłq��\��g��9�O�)����z�`�#l���݊�6 n���S�l�6'��hK�N�ky���������J��B�=�	�����آV� ��H�<u鬂E��4���ss����PRv���b��]!!{jr̺Sc�cGp��t���z|�Ȉ�vW
F/Q��`