XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0%M'V���E�bt��x$\|����=���3�H����m��n	~��D�:q��u��`��a�e�C=��232�P�
��q�,�t��� �_��{㐙�3fk��J X���`�"]�ش�Ǒ)�w�O�������Y�K>Q6��M����l\��kK)*�Pg��FC��F{������'"9�KJ+����Q�t^�7���/�#cK:�0������Q�'����f�w�]ks���'@+�i����=�ףA)��ĕ���U��T}�61&����(pm5�Z��fu�C���U.Տ7d�~�)��t_�C��4���0�V�7
y�{"J�g���T�N��B��i<42�h�?C��|�Q濫	������G���E�J[�߲I���Ɔ9�Cz���Q��y�|ѠLs�'�gI�'�׻�<������xz�D�!{6��ZL���v�OL�)��m��(�a�V��{Fρgce����3�Tq%�2@�����Ϯ���y��T�Yэ��(Ϡ� �#��H�-WxI��zsUwi��t�X�T �y	�^+Bf��l�����N�h͘�"e����^q e�FNl=��	��[^�@]�'�w�䑦zUw�M;ɸs������]?��9t��L$gEr����6E\(a�w�?SӀ��� e��\K;���-���k@�B����鯡�(O
>5��dOc�[b�*|��vlr���̇:�=�Ha ��'��9�{�,�k��ܗuQI�XlxVHYEB    95d3    18d0����4ۘ�J��Ϊ��m��n�1�"
{������0��%_%:;���Y���ቅ<��fz��[2?�Ķ��7�IJ��Ⱥ���?�O���?��lv6 DF[�zv 4q�`C�G��
�Ǿ�멞�;�P/{v��ޞ1��D��_A�1^dH��Сq���a� &Iu�Cm��c���;�m�nN���"`)��^a]�����P��;}DD�p�F�I��Z�.�Yo�f	���ǜ�t7V�HY��kX�Ú�:����UL���0��E!��Ycʎ"��2<Ԋ�����R���R����Ţ!��7�|eJК>����GAjO�g��K��:nz�ĭ���/�m6��aO��q&��ܐ�O`et�Z���<�Ai�P^sBEs�?[��' n��/AIt����N���ZLz��w�e�y������n5�|�./�|g��,Ʋ1W��0�g�d=��0��g�	�#����@D�1,E$�$F���Ƕљl�Wރ� ��+ds��j�ѷ_T;�"U%C����O��)|��z�w�BCN��O�*��ERz
@�`��I{a��6+�ﰕ�C
	�q�n{f�j�v8�#�� hCƀ'%>%��<��W:z�~J��?��_���z6��1䴧W%�d��v��a�Z�]"ܓ�4���凤na�ܰ��8ZAi�� 5�^i�[|��8?^rC+\�]�Pz�g\���=P������ݼ<�w���R�J��W���Կ|��G�!15h�!�:z��4����I�9�s{?|�B���ac|;��9p�
f[�V�����ￊ��&�_j����2L�]�	O!���˨�ʛH�v��T<���K���[���kR&�.�r�4ֿN�@�U��~�Uo`qs|������G�{'F�Q� ��r���R��Ni�b�9uF�U*�eF�m�To*o��k��0��	�d�LL���2�E?�'�-dC ���}�ET#��������{Y���o�����2�*�߽���}q�2T8����oK�X�|V��?����O�q�V,��7�Y�0o�X^�X��Ѧ��ߟ��j}���!q.�GЊQ�����4oC7��L�X��D��l�ʋ>xe���H�MLO7����k�!�B���C�92�����#�w���3�a�T�%={�Ӡ�B�[���mv�rW�4̎`JW3��h�c�O��~��>�Y�܋���
n�n�F��nia��GI;�x�&�_��W�G�4��t	
��p�gPE�f�Thh�ܸ8�j'>`X-|���O��V�}���*]�߄z�&�H�u �r	�^U���qp�����>#dk]"��o�8FL������)�ྌז�Wz��wg�ajC�'��(�=h��;����y�X}��_�]��;C�o�Ɋt=pl���'#u��󏜃)��U8���zt��W�6�D����9�@�/�Fz���W�n�^V��3p!ǭl���l9m	�+u#x��p��(�kolk���fs�O�`Ƿ�d:3���j_�xʈ���iE
�#��U��o��T�N����V]�T�ƙ	I�Vr��u�I3��v�0��5�L�M�A��x�'0� �phV(9�5D_�xȆ?�3N��Y�����R������+���[��!e�Q���N�h7�e+����:j���[�� ��3���dxe.��e��2�y�Y���j���甐��Z��eh.Al'F�) R��ȓ�l��	�\�K�����y������%[o	�g����O������kL9Lh/�H��z�EG ����Wi�e��/h�~����A��/���\��88�:����W�\����L���v46��X��U�8|ԇ��<����w-��GGўIR�~=�bá]�Y���x
s�`�V!��R�LҠ�"��L�`��-�(�h	%���[�8�pw�Z��d�c�:}�0k�/��#2�9�𭬐�̛0�a{T_Jрa�m����;}^.�Ҕ��>�Ξ��սw�}�w�� ���OT��m�|ގm\��걞�n�?����ycǣ��Ňn'�ݞ��S'����ӌ��[���݂Rįy5��ޡ���ߋ2�8u[8,}�p:�o� ��	�`��4��ejC�m�dR�mnC��Ӥ�z �~!~�.]�^����k_06�[�_��] ŧV��5��/_i��br�2�*3�0�+�?�o��������F7J<[���B���	��L.gvtvϠW��G2$D$B�c,��>�����w��d��.]�y��̞-H[1U� b>l����?��2�]9�y��O��{��;dҰD����(���V���kcy"f����BN��*m������K-�E"���iK��q���+wJD���U	��HC�����i�!R b�f�\�r�>S`���8*S^��-��'C�E����0��c�F�O����r:�
@����5�\��V�[��67�ɇ.y��ٞԦ=`V-��uES���� V:�Q���~T�I�]Y�d�k�M�=V�!������3X���� �>��Nqv�W~>�ܓ�����s�z�S�ŁNi�4�Y��v�!�[���0�agg*���|��@	=�����k%���._n� �;N�����Y�Y)	�r���56a�J�\vv˂A�A�)�B��'�k�e���T�z�-��4�cVM�w�ec����),<l��[�D&�gE?�P<��&<P���ދ�����B���f�N	"�����/�%5��t����h����h^���"��Z�+�\�{v��%O�.�|��EZ�a{���V޸`�Jl�./������&���+Y��C�f��>o�,Ӳ��5�uJ���Ǡ��3��+�H��:����u�qXl��JNƝ�C�-�Kp�N�� !P�>�5��6^;~K�Dw��ҘPU��@��ֈ���=���.9Ls�<�+@޼��7]��IMz�F3ݦ����L WO�y�,8z8WN�wѡ�9��p�}�$�Z�{��� �A����*�mv��Uݶ1�*�f ��}l�8=Ee^��5�,�����<
ܯ������J̀��k�[?���[c$��ݳ��r���/�çf�n{Aˤ^�� �|�����'E�����U�|6�I��SZ���,�.�ʑ\����ɛ=)δ�=�aXb�?:몔�c&I!��@���7�-��w��"^��f�OB*%�`S<�"D拝�������;)-�\����m_�S���5K�q�ǅ��~������	�vC΅m�'E*�?�yf���g�Soe�C%	mͩU���cJ�#�.��<ո]��*�*Y$�Aa�7���6�w_
�Px�;�|���
�u�ؽ���&o�k�r稆������������C~V'uG#�6�5</Yʦ ����uI���'���NT6,���7Ch����؜�-��K�&k�}<��U
2_`F}x�hQ�E�r� �V.^d����րjי���xZ"����վH6 ��ƨ\��eT5�ږզԚs-����FĔ��YA:tY�嵻W�������o讦G6nP�u�%�"���G+`�S~�	v#�S���-�!���΂f	ye�~6E#��)m(6�W��J�чC	�e�|]݋��ey	�v9�|dx���:�r���p6������]��R=DA	/��3~!v,��Ĵ7��G�8Fw�r11#y�N�	��:.��P[j �2zL���[�tק�$o��rƒ}`�,1{�~f��5�\J;f����=� �8�5����|�[���M(���{d�Kg��7s��q�
T�Ce|�k�}-��M��{U��,HʥN&��6�X�	���^G����|��&�DK�i��w��r�G��E+�M�p<K����iA��9?�!�tW�Z�n�V�kз&`xU�X�;4B��2���}�?����}���C�s;�^�P�/�/���~�����'��z�??���؉<G4�{�+o�����|���������Rc/�WOn{F?������-bΜ9����c�����`�'��R+�+s��*:R�Y����&Y�wk>�2��h-]}��%o�GT:��l�#H�u��s�Ճҟ���9�Wd�g:�_4�I�G;�8����^��k��Y����~&������68��*2�Cc��h�'(Y�ތ��n:�	bM�,�������TÐ5ό�%�j$Y�����хhDG�ŉ|�N\
3������{��<��MQ͕X�R�u��IA�y��i�"��|:@�S׷P����t��8�p0��=����:Pk�ܰ������u�q���oh���H�H��	�'�.����う�G��L����6*E^0�Ǩ��2���z�.��i�cpt)R�7ݖ��sηחJ�`L#}�¸�EC~ʿ���a�c"��Q�d-� �VYF�����G�S���w���ݸ.�JЩH�����Y��	�l[a�g�UK|w�\å���V���+���v��S�򛖁�竎.;{�^���v�١2dX��7�J��@����(�ь4��:Vڹ �`B蹋��Yx�n[�f�c��K@��X�H=��zj$���l�ia�i�����B�sX�\M��6��a�x��	�f����nbK��%�B*_�ܣ��ą�C'#X)��Z�oO�.E.���`r����j\	��u1��<��"�۴W@�?������DZ����	 fp�
��>��@ټ�eR����=�������M�~g��|VӠ���p�8����Ei[SʭV#��5찏�Y�?l�����!%���������3u����b��Zǳ��Qfl�*���5mΙo����Vˮ��Kg��|VL�ΰdMz�)�"��TQu9f��?-g?�Q�CP9΅NVr���Hx[qK�?������.|�u��0��:��	�����_
��|������� ��J�X�J��B�7�ќ������_�z'�5^�kj"��f5c@�{��x&j��X��>�@#��n��sH�1�|��,̐K(6�eU��OX�>���w�]a�4G�����ә��>%�='�ieM��H��j·R�8\����>��G��y�I��k�~�5ɀ(}���όF�K�nl����@C� �n�6���1�8�w�=�SG��0�8�#Mq�YBc��$����x��{���)DFHGi��MP�F{d�	9ME��c�%��[.�&c���>t3{q옊�����?u� <��&���>b4���o�'�̀;�u�}����y�،�K�^�O�Q�1����� S�I��*�n��)�6����>����s�:�y�����N	�\��5|���	��>�l9�����T�ᠥg/�8��3�}]�����f��cl�*�9�e2lS��ّ^��+�bh�JYE�`��|��8����R�t�V|�^���B!�H�z�G�e���U:�x�|�*�أ��kX�(<Vdk�\Q,�Wų�)X��aШ2��]��_2`3�AGɮ�Ų�sMd�]\�x`�gV1|7�j��"�\o���\���"$����n��k�NW�o&�"
!�7i��Bk��1A���c�� �Y���H���B/,=g�3��:2�F�*/�(�ǗI��^.U4v&�ҋ�G��M\����@�Eu�\ 2���K�z���Ö%�f�{�H���i�8���:B<=�ٜr
o�Q��$_y��fT��=��ě=,Tߺi)f܍\�:髥�>����Z�9��Y�%&ش�meN������ӽ��rMO[Ta�;J��� ��W�p��3+�-h��a͂��g��v��u�����B��PE�ӝ�C��n��ZտG�����O�~���˕����.����[������YX@�/��j%�����&	A��1)�N}>T��k�¸����*�0Wh���u�`Cϑ�k�*�G��W�����Kj+��3�V�%jZ(C��&�uܚ�-_ ���?���6��F����2�
�5qJ �1F�]�����Μ4�F�e���y��ܠ�Ey���&O�_��6�\���#��Z_ۏ�ɮUP�@� ���[^���A�$�T}Fkh�����W}/��rX��>,�o�� �JAɒ;ma�b���mt�-�N