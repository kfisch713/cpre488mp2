XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Ui�Ԅ�V��G���2n���pb]��IJ���-�%4IY����[�p�}��f�z{��lZ�XW����d��	�������v����t0�u:�'�_���������'���;ݑ��g���ﰔLZb9�5N[�`�_�{�6g����K��?O��䚣N{i�O�����x��b^�{��93pv�,cN:ٖ3�'��~���E˽e6Nl�p���n�>��:t���`�����������b�nX��*�z�0߹P\"���,]m���DZxQ�:�?�Hi��|�Re����%���P>��-��� O��1!����&!{V�(��Yd���צ�z2�bxtL��K,`�Z�D�I�^�ѩ�����V��6H2��Zq#[����43��Ԩ�OY�5Ix�c�|22m���G+e��O�c���L� ���n���+��qk0M/��c4�8��&�*[��}�[?+�ˉ 	]���#�x����<�����������N��	<���m#@�"쐢�"�Ȗ[Q�z��	��/w�}�/%[���=��G{�D0cT�A�2�;D:1Y�[����
fKRH{�	�(�P\,�)J��r�#X2+�5sjML�G������<�<[��g.�4_�WS�ԧ�]��Q��4�ɛ�� �8�K�v[��=?����tv���Ryv���Ju��ȏ�&�m��>��P����r�5����3���\r.c�,�-�<ҜR�\%�r�i��:W?[��Hb���XlxVHYEB     e07     680G�.#�F(Gf���KoE��|{��D"-��O��k�>q�U���m�>�S�UE%IϏre5)'���Xs]4�=�=h-֎q���[���m��aop.qD�y���,Oq|���L
Ѐm'̞o���p�١�T�wx���`Qt��Yã�ґ@��H�(�<�<�,�(�U���������o��k%���Z��+�����&yT˳;���Oۗ���t���H�*��)��Q,�|�[j�CVj�@�H����u���� �#f�i����ڌn�-�*/�QI�i�zr�ᨸ1["/��^w���H�&`!� Os��yR���Pr��hOu��>S3-�drXʔk�|80 ��J1���)�8�XA�23�̫��/#w.�ߺ��I��j���������P£����U�߷:�o���<��{�ǧ��Ԥ>���Ԅ8h��8�+y�{��l;	/\I��K[7TŐ���<� �)!���.�hW� ,��L�<�ivϺh���\��ݙ�Dt����/��f�1E�\;�֌�Dq+i�U�1�[��?��ְ�!E�w���V�mv�P>�Y2Ŋ1�Nݰ��%��L薛f��K �h�Y٥��>m�>��u	~��7�,��V.{:�Ubn�o!祺��׃78����ҸOb2�3�Z[����$U��Ua/,`�݂��.�
H������G�����@y��7��(�(jP��^_�
���_`H����dO����/H�ci|�r�.I�oE67�L$<����Y�6�f?�B�$���1c_�f�u�o�;���j˅�q�y�`�i:�����v�}Nؑ�S�����r��
�kʯ��tY x�q�(ՌC]�\/U������"��\�DGqO֬���^A4o�F���L������s����*~}f`?@|�j�H�u,��X��� 56����fN������n�s�E��X◎��"w���sd47v��1qEs�X�m�
�����(���5\��{��Y
���^�G��z�:�P��4��:Ҕ@O��z%�G�8��d��պP�;�a��hZwՃu�ln�����FԶ��B*����ඓ�&� C؇��;2-�(Fc������f|Vy�y6�,����	�-vd��ڦS%�`#�o$F���lb}��9�m!3�]�b��1U���3R�#w�l������e�u��
>Y쒴r�[}�O��I��sm��"b�luA8�����&{j��*9�M�[�r|'s��ǔ�X�)7L�)m	�W�ur�c�=�YI��(f���1��D�aL��%�\|�#aPN��F��d�\��������U���_�]�PFXBv�:,?����2��ͬ��B��j8�X6���rX;U�|�Cق���D�6�)��n`�Еӕy�6U������F���ëk�_H	� lH=��/�j�]y�y,%ؓd�`[Е���6����b��uMz���ݿ\�2��� 3\�WC��N@RHU?�Ú/��(�)�7s�M	�D���<��N����R1�)�� ��%��R��u9n�6�>������S3ΰ&j�>�\]�05���^{���5~�U��Q�S�Ҩfy�`���@y