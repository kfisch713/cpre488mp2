XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���YMbM��]Q�����
I��H�8��M�ު��3�Aj�B���� �#4����S?�{p` �NpT�#�=����O�i~+���swD_��H&7$����d�֎#8��+ft�i�	�vږ4�'���v�p1��QrW�U�HV�x�r���M��-�J��i�]�qONvY�*S�?b�@�D�p���9t���V�V���F������iJ¶��;��h!F�hGm���0p����(���O��߯��p������1F����<��g���a�pu��x��γ\�9^�&T�n��/Ck�y�dj�vi �:[OѾ�[b�.�#��-?�(E���
,y�Ii��Qŏ>���(k3�[�)m�\���}����<'���Lz6�,�U���F�}��i]՗�=9���|N�Vx�3k��f�àq�OZ����{G��zl�I+J���f"�-��.r�jk���I7 ���`��ӊ��{�G�+��Ձ�S��ap(� ���� 
�8����z�O�$"�t��왆� }S��N��$�eoL���G&�yь�<B�5f1���+?Xx�Qw6��и ?�-�rL����\�����q%#��r}��W�5dZ�!�H��)������{l5�_3�Z+��D�6�E�V]�%P��b"~(�Q4×8��{���CD�i8ؒ�����G��%�,N���1�7n�[K.�rD�3*|]qd)��^�oxKs8��n?{B��ҏ��ESaA�dOSP�q�[�z1�?o�XlxVHYEB    2892     bc0&��'녕5ښf4���,v���wT�� q��`��8��;p��s;�xY�C0&/-�� o���o�A 	i���F\HkC�e6�v�jg��8Ap�K�����CܴB;�u��(��(��Ƭ����@�</��MӌX�PU�2�ufU�"�5���r�Ҏ%�`ʢ��ͨw����b$�[���q��`Oql��-�H���Hʜ�p�JwX�W0"T�6����a~�%u���|��"k�v���T������
��6Ha�m�Y>5�;�duTbN���F���e����>�;�a8 �L÷H����vq�B9�-\D�5�Yj����@�f��&Xd#U�'A�/����.= *0|�Ӷ��.��6�8@O�0���z`Vt^��JDO���� 1|��)�H���|��a޵�?�k�Hu���ݏ��B[�z�@��bH�y�	1*�X��E���8�wׄS��b�M����X�I��l�4G�o�!
���i �V��M%��V�K?F[��r�e���ׯ<��ߟĳ��/�F�,2ɞ8s&P��ό�������4�rV�W���F�P�."t��?��U�2���<!�y�m1��R_i}��8xo��3�џS�������d�?at��F�{Z����	�8%���"�p`Td�i{�^�}e,��UH�c/3�S	b�H���I���V����C��l�T���4�c�`�7�mJlKu���V*�W~y��� ����2\K�'P�M�G'^G�g��n�����T�,�w�����������&�!�0��s���n~��骨3��àE7Mgf����=.�Mr��Ė�y�~Q ����'l�qE�w�cP�q�
���
������J�9
�������|8��n���eJ��JG�2��ɹ� �?i����9��~�����/1U>��kG�О�lk��ʐ�泊�C϶o��󍥕���ZR�|�Nt&׮�X`w��˶��˜E�-�f�1��r�v7�e+���Q�dO�J�o.|��ub�S0�}���1Y.�	0���j!ǿ�81ΗM�]�3���<�)l�t���2C�(�Z��E�����5�_�Ce/Dh�r�7��x�O�
/�b+C"kg\M2�-�$��4�(�"�	��pp@~�����6���K��u4r�&�,+�uu���)� �g�7���PsJ��Hh0��GM��ǂ⏼��R��=%�q\�H�>ljsݒ�"��ͺ\�BM�G�U��`��O'p������"B������2�b%H$W��'�%#י?J���Ū��~�$GL߄��Y]>��W�(2!Ef�+�	���5kr���_�{Ex0���X��A.��pR:�~�^u��9��f���/*�=�i/���k.�|VaR��!�?�a����R���'��'{��k�X5�:G��"�(Hs�7������VM�cu�"V.��E��'�Y2@o{n�L�A4�a����R^��ʬ:2�s5T�v�p�c�T��x�k��r�űe��������G��&���7X��#	�H��*�Ϛ�N˓�.>�X�qD�5 ��6Z�����U��%*M������I��x+�Pj�b7��+�ܻ�uj�p�`��%�����RQ�<�榣�QwD뿤�樆v4+�C�u�������LKڻ��Khskp��	E��3n��G��+ͣ��G��?�{d���m)8�<�ɾ8R��j�)[��&����i��6���R,�cJD����E�Ul��4TGx*{����W:{*U�i�s�N1㝥P'v��E)m���}�P ��fX���;M����jH@�>��i���I[�*(׮���F�Q�	���~)�<ւ�}O�2[�8�s�$��#�f����ʇ�7u�k�׈�l�V��i����#�7���@/F{��|��*���M�o�!,��Y#M�w)§R�Z����?_Ѫ�<ኯo�\�K�Ս�ʬ��=��F�/[�Uf��F���v9'�ֹ)�OU=>$Q�:^	�b���q&�j�%�Ǚn`B����ZC�G�����!	ĸT^��]�身��d��1�X�tnX���;`�����n^���E5r�����e�<w~7ٱ�����ds���k8�!��;��G�o���[�.=A�q�FM��ڿ�#��+}>�L�@�q�"eu].�8s�}����b���(����-%pF>��Q��{�����2$H�#�Mc$x֥O���=FUsm��Y}^��q8@n�[��ᅒ�<
&�#�no�@�� :�m>��zI��ʌ�ŘNh�{Rd*\���4��_6�Fvw�ɷ��:��q�=���V�]C`��m�5:I�	���c4Л��44����^�5-�٢t���`�g$��jN3m��̵��D龉�T�c�'ͦrgw�g���9�'Oy_OOb*чZx�;D	70�	KE?`��Ʊ��%9��s[@y�����)RXрP��b\��1;Yaw/��h<T��z~X�=^���¤5*4+r���i��ZtiO3=(�=ȼM,�	X�� �W���Lw���N�\8�b
�,�a�ܣ�O�n8����-��[T~0�i���s։/ms*w��("nAٲ�!���Ju֯�9\매9=K�")�	�pd%U�]��H��.�D�H�85����H����h���iTg��~H�nz�62"��Xڐ;�vM�ᆄ��u���(�lv��eyb�=V�dt1Z���6l�E�$�s�s��/yb�o���R\���^����/:�7h�Fw[�������G��)Ud-��N�"J/�O�G�t6eZ@F���8��%���	}m�8��%&b����K'h�n��b�S^,P��
���z���y�Oa@�asb>�4Ȭv73n1��������rv�d��A�4���v"u$���U0�<�?n6ol͈x�g:;#��