XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+Wo{�^�vԏ�|�slWY"�+1�/:�7��z��|~1j��k��v�H���H�텟;p�*O�q�hD� 0,LR���PQR,
o
-�V: � ��/�A_$�_D�u�E+�=�׶C��8�DWO?�B�� �[C��
�L�PR����ň3ʽ&���^���fj�� @��QYIxpjY'ڽ'�4Ɯs�TX|�Q�d'yq
使�"WjY����g���]GCz�򍼑go(��`D��	��ֱ�있P ��A;u����2D�[��Ӝ�T�|��މ���9x���0H�5����4�ϔ(HbN��U��Dm��!�n��}����u͏��Л��������~�}���)�Wn���i�|�B��_�_bDR@�.��O�h���ߣ�M��C)޻�:����?���Q�6��n��א���H�gݱ��;�3mj�we:��N������I;=����(R_+�'@	�	�9�2L{- B��%14�"e`������dX�$�j�ͱ����$�|�]$}*-���g����ǃ04Ԏ�n��������qGƺA��!�<6�\�26aZ��5����h7�㽊(�x '�����,��lݞ� �hۧX����b�=z����C�9u�D�n6�T%�9�]_�r���S�Eq����^S j(إk\�p_r�t�7��q4�V���ԡ��>�_Y�l
3�emV�e�J�dV �Q�CP�T��2=�}$�4e�1jT���!D�����_��]b@�XlxVHYEB    48e3     e001��+<�2DC�}�G�F�N�[�� ��E{��.��.���l�[�6Bn>��<�G�5Q	��G���t�#m��ک�1ê��y����&�C��T.�"��䯢0�)�� vчQ*#�4Yu��$�m�U��ilMI�ښ]�L���M��N���цڸK���(k�Bs�ޗ�9*��P�DB��F�m�'��͐t�r�6�>>�n�(�E�٫�VB�1$NWP����T�`�9���#}k�`��k���`�9(;>\�~���f����z�u)�o=�Ŧj)�$�v�B��lGքs��4�5��S _�e?�*��c,(^ČM�7N�JW^��[ɫމ՞��I��.�r���G���C�'qZ֞0O��c/� P��!)�!#�_ ����r�0�����:��-VL1�uun%<�n�7�Ee%���E�,x���mF)��T>�s�l�%n�46��%+�p����ȉ�VX�[����\�a�3�Cx"ќ�];���xI_b6�e�<�4�|��¬�m�tՓ�`�[�,�Eu��7�'� McЈʎ#�+���<�j02E.���^�$l:�a*:�y�C�Q��n��A�=4���*���ܐ�r|�5E@6�z�ɵO��O6��^��\#�c�g=�ǘ���ʄ��
ͪ����;�Δ)ٹ#2���Dʮ*�8�uk������@:άX�,�tX,�����ܻؼ�j+_�W�:�
� ��NĎ%�Y���s�w����l��H�Rpx���:������!�C�o�H�h��,�e5���A�I��w�+9���Y�I�t	���su2_J�~�=?�7�ہͭY��R1����X�������s�g�M�T�;H�ܠr��{q0�6���.�S�E�w��VP.:�K���gyD�l�5����,'�8��C �U\��E!\ƹb{p�Bz�u e��ilڻ��nD·jܟ^,�y�G��ʜG����1��(��'<�yۇO��`��0X\�E�o54�_i�3��""\ �K׼O��c��ɷO�뇭%i��>�j̅���f@u�M� ȼ��Th <�F��{gu!�j���dl�14וa������?�ۛ����he�����GVa��;������Л]�k(�.��<��O@M�2�ZjIz�[+x.!�� InGwq��B�B���:`����VD�%W��^�,B\��U2b��h��e��x�cK�?��V��H�ln"��!��g�r���9O��wp�%E�Lz^��ߎ�(Z��Hr��GT���젟а\��:���s�;����D�n�U�ld�-X��/4ۆIdp͒��I�H�ʊKy�2,�lu�
��FX8ܗ�e��Y�i������W$²~���؃XG�T��])g���rq~�o-EWqof�FŖ��5T3ݣGd���l�G�(*Z2�	X��H'�v��qQz��zY�l=i�-�<��������*�9��y��`��*�����A/,?[��n��q�@�Y,WC>��uu#�|��[�W�����:P��q�h�؂K�zokj$��L��敳�{�R��qK�v6)��FE@����H���0��;Z��(�M��Aͷ��l�nf�Z�/��ߠ�>����̮�����Ⲧ�נi���u�r�m]Բ2E,�o�/y�Dk>�%��>:��/֣E����ng�os���T��m����,�qѬ]���!6x
w�!�^�������&J1t��g�D�ސL/��Dy��6��-_�>rKjՠ�\--�1��s},R.2�UD�;E��*Ia�U!B��7�d9����o$ˇ������ ����A��sgk��Ӷ=\��zZ(&�p���� K˦�nh4��("ex�<���n'��e6��	P7��T��x��ĥ,lm��w��"1�"b_�,�� �q@���#��D�)��W}�|O�nށ�Y��puQR�KlaÂ	�욤#=vKOXiMp�ry��O&�xA)YtPd@������5,�>e1�V����/���i�� *���$p� ����2��)�p�)�n��U��ev"��]�);��'�m���ת�9i��N �IϰY՛��z���go�V˱���}�9���'���}khۺr���qk�E2�)�i"�"��vx�淃��ZC��rdu�B -F����Ө֒��#uz$�B3ỏ�y���y^:!6���u�"Ey��O�d��G�bZ��p�A&��j�g�����e|[|�R�T�2�7&`�����Nv'f��MG}����}(���ɫoc\�ݞ,!"��$��<��⺇���&�3���ʳ�o��0G�+�jLIg�e����s��ˎ=�lr��c=��D� �ϋwv�<�HrRi\Z���66�|P�gv����\���-ݕ$��= 5UP��Ut�&��Փ���ǬͶ���@@4a~�ޟk���*�������i�W���A(
���eg��q��KC��`�y8Pf��d;��0�A���¶%�/��Z�3�L�\��Ϋr����c�ңC�_?����D��P>2��w$��X�0S/-v=�( ����0'�(Х�`�6 Nf~�i�8 jR`A��<�n���8N�U�A��M���/�#/� r��V���VL�հFN9�i�fߟG�%z'yv���P9��Z�'��'!Q훕=���Ɂg�����0���2d^�[��>k^ྏ���O������}�Q���7�3�$��� �U�yc��:��%3qT+iu��t�ͷ�����pa-���u�j2���;�Fτ&r���%�����P�������\�KG�Z7�L�׸oɋwI.���tV�ե���[Ǭ61p������������$�{؆FE�#�i�Axo�߬�G���g苅"'r��X��^'S�+�q�Q̲�z̡�����v{���uv=-po�S�-K�Qw�۹ƛ��K+�_]zA�����u�}�%<Vϓ���f��s��~#Rމ�YZ�:�Ý[J R<�e����5Y��DR7[4�LJJ�� �[�J��}����x'.( _P�v����[�F���M1p����u����	.��0RW٧Q���#����Z`h�;�$ޮWBb�4{�q�|��~����As�n�uّ����������'��:bM��d0��s}�\߮[�]w�1��unwW<F����5�B�!�A�?9�/X��耇�i�G8�+�e�xq��D�n���?���
�y)x[��Ǚ�;o�����T��͉*��-Qϼ��d� 5Rx�}O1m��ND�4�p�$��U��U�Z�� ��G��W�|@N#����_W��bjey�e��t+k�h*���,2б-�{��+0�qD;9��E5];����_�f����v��DB*����
�S�ws/� D(�?�e$&|~]S8�9>a�Cm�Gz�p�!�w��eWs�����o������֬�u'���� 5Dk!��6|F�G�H