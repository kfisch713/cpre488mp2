XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!Z���tz��~t*���H8�NW��$����I�1�>GBFh�BH��	�������Z�}r�"ϤE�M8��G�-�iƷ����I�'�[?�}��������P���*�+�\::�+��9�ި�~�x�饱�:I�^@�"����~G_�U�So�Bdi�U�&%o"��<isG����Ϣ��ړ�+��?�Vh���I3^�v�]]�^kW7RL�8�{�����;2��>0���'Q��5\Vja
Q:ɾ *�BM�d7Ӥ@ȡ_��S�711�O�2�KH�3�4��$X�����/�-o���'t��KEM��^D�r���<���o8t7��cY���u~�.�7o�݋���6��{�2������g �ܻ����I�:����:�s��h]�la?H��
m^9�~��ā�ـNd�M�����`g�渄L�٢��U�r�J�s�9z���%L���&^=ҏ\Z�g���Ҝ�H�Ѿ���/�-":;nO
H���FqU��')��|��+i�1��XvdE
er�Zm�sٺ���؁k���V5�]� =�2��PS��#]˜	B�~� �D�~"�a��޵�4��6L���E��!~�F�~I���bֈ����
�Y��]B~C��k�'͛��U�'�3���]Ħw��G��=8𠜶�C�GY34x��_��@�n(��W �e�+ڥ7�Օ]qF���y��=`�G��)��g�<s�~Rn�h��^�"w�(/�*vH����XlxVHYEB    17d8     890u����CA�1	�A%eJ��A�^�	z�o��MR�"��[��M�UqQ�D'iof36K���0<c� d��d4��#w���z٨Ci��jX�Cawwp�&;|��Z�L�\X����r�F��Y�V��կ��9�t�*��ީ��>$:����5��lm��j�j��Ʀm����w~+`�h#� ��?�T�Z?���
M�̎�����$�0K*����G����6Y�l�h��H��N�#Kk׹��m05���i$#��_.JC�mM�O�F_&/�JG��i�x�x�b�1�}@�t-�Y�-V���r&TZt�EhY}�vF,���{�g���	<�����Y�m������1@DM��j}�r&��i����V��d��3���5�����tow�(��[�L�XX'R�}Cy���d�EKRߗU�"��B�b1���l���-={Д=1�]\Lj^I��wֲ�z�Wp��f4wQEp�d��$���
D��R��@�;�YQ�s	�(4mZ��,�$I�m�0h��#����y܄����Q+8e!CS���2�����H'�?5�J~A�
�l��,�ZC&sFsSl��2?�<�O3؀+�����s�J�+�)n3w����v�h�@��?��|U��[!÷��)���fC�F���&������/�WO�Sx{L�j��:��kg���b(}m-XĺΠ�k��%�i�s��_��N�{32�Va~\@x�	/��N@�&���:N�]�Y�T:�Y�>H��}w�r�5�o�,��j�k_�4��7�Ȯ�+E��|��-��ؓ�&� �J��<y]:���~�5�_�s\韈hK�l>�6�m�;�CL���ax龧�=�KM�[�שgoO%��]s�?��y,"y$>U_�����Y��c4E�\%E�[F���!`����޿�5,�
��	����8�b��*�� D�;t!�k�RgG1�U���+%<n��jp4)a⅟�R�6�kim����]����rv�9��*h���5.l���)N��)����ml/fMl��%s,��KD�
��ɼ]x75I-�3X�����r���gkm�O��c�O�r"�9��_o�����j�p�ҿj_�3:5(��bG:���.�>�P��K&JѮ\vӑd��餜�,�C�\@�"�d�&}�U��L�j;q�f�!�}aB\������?ۖ]��?4��%M&wh�e�m�,
�\���Js��I?~����J�8�ӹo�ԃ�|�6����՝�3$�%Ր������Y��U��t6KA�nxH2�oQ���u��Ħ�6jh�ՖR��h%���^W���֔vm/N�?$ꭉ��QW�|2��T��C�*p��t�iL���o�f�<���tLw��+�n�;Q������F��$%�\^���6?�ஐ��@���t�A��y�8ΖQd���g���@�6��ڵ�۞�-W7h-���d����v-V���q�OB�Y{�S0Wq��r5�X��o� �z��=��e�Q��G�M1���5@><��"�R�©�d��"��̗���*�А4^��,�`t�"D^xa��;���'����
ܥ����:
i`���4u���2��8�L�l�^�)tp�ׯ2����଩W�lv�3q�~	�x�8�Û�c���=l���\�_hZl�g����č�0�=^����'W&��ŉ��Z�#��p}��Kefh��f��5����g�W}��Z�OM4�W��l��&����<5�����۫gJ�y�� ~����b=At�[�;�t 'k�+��gi�cJ�-4d.�����*C��w\�vuY����HCt���.�U�>уWfӼ��b�/d�c�&�p��K])���P�1y}h=M"������#
�e�zp.��=.<�=>��ʹJ�z�2�93Ư���ʩ`���x����7���:���jXL��8���| �QK�����Ye�3(:�w�5?�"!�!N�]�Kc����0\��&�89�|�Z��t�@��Y�LL�,�0XN���Sk�=�8��c��nQ[P����,M�kS8��H�m��Ս�=��d��x/<��T��P�YCN1E�۵��wn���P+J�W�lc�X�Q\J�����a����*K�*\�p�