XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:�������B�r\�)�KSR$���B�m��U�1�_�(U^�Bu1�>��ZIe�b�TT��ߪ\wY�s���M��&���S���8K�g�-f�X��>�r��H�)V+��Y��VZ���=����4�J��>��"
%o�B��O2E���./�}�Y�V����s��`4��Hw�$eTکU�tk?O�3:踢'+��mG��~�����Y���/UZ4q��aF�[݅.CbZ���d�z;`�)�I&u�V�@7�<�ck��sٲ�\I�G��J�*�ײ3��sN/RS�&���K�s�l'�
A�.�Z��
}]/�^�k��I��m	�A�cU�>'��IrǼ�곈�ۇ�eaev��=�z�F�iG�����9��r׮�:�NpG2�����đ1|��^n`2up���Qԧ���L"������Ӂ�]0�jr[�M��?������]����S�VL�Xow�	(��H7c�����0h�pJy�J��N���������x���h�q�Ғ	'��o�����P�����J�Z`ak�%��9��-.�,c��������Tiͺ�<�-�W���Q��r�Ur0�j�j&��Mr�䑜��ƈr���ycg���_���p!�K�����9�EH��+�5�b������z�[����F(�(�6�+#E~����p��.�+p �;vl�e�[v���:��=�8���Z�����4�Mq�_�7�^�JĿ�i#h���xXlxVHYEB    3fdc    1160C8�3���`�C�/�v?[�;�K�%2�g��Bn�.6O�rF_�ui��?�0�_XXj1(���-�,�;�J	��`����2жMtJ��H�3����ɖ��d�Ceg�*�����x��K��Jo१M�c�����Q��v��c�t�\�^7mee��t��ZU&�2,�қWdcP��Q�6�O��v��`��X��1��PrӚ"�K,C��X΍l�:�=F=�є�wZd��Vk�me��-/GY�tE�+
�_#aB"�^0�#�ݸ�v,>���� =��ܗ556�H~i�$���Ng�'�2���BBf��o�����gqQ��	���!9B/����a�5v�IY�p��l	3}4"��\���~btD,��C$�������W�ǻ��#�e��p�H�wQ��t�;�j�i�4>�Y{����K3�B���u!�c���5i�+�v�}o����ɒx��G	��<��? Sߓ��s�L�}?U!}J��'��𩼠ʗ��kˊݭH�4!�=��[^��dDw�=�Y����|�v�RD��X(��ع�Ǖ�C�<�?GZ&quď\� �z�s��r��ـ�;�ۥ�Rȝ�SU
3��3� ���F.P<�^�j%$l��\�&�qE9�8��,���;��7%��G}+��'��ò��c�� �B	�3���� �؝(��&��U����bs��=��k��5\�H�zW����d�[���M���cF��."�?��H�Cs��KPF}< 9i3�"b�2�3��m0,�ʴ0#��	�M;��3\]�	C��A/�ʫ�4�DB�I9-I�\[�l�F:�|7%>�s�N0���]�d�������	�}L�B���lxtk�B�Lan�'❌f��4Ծq������R�����wb�]� �q�)�n�(�'R���k_D��"��&����.��z��t<o�3%�|	@��c��{?��,�5���*ا� �t�|�H������?UOY6ɒ,��;����&
�Vv�[�e�, h��4x��f�>X��̀$aկyZ�5�B��C@תu�ar��v.�i�=ב� a\[s�^H`��;�\��^�i��E�-�*P�1p�o��H"�N��j#DV��T��Mڧ��E[���ĹX�,**tk�d0P��nyF�/ሂ�v`�MT��m���8�E�&	�q<��}�/X�C���.�E(������/��	Ζ����VE^�]Z�#��3\�Z�0*s0�x��u�'X���u��Q����h�úAJ� �|��M�0�"�3�uф����B�@Է��Q��Wȝ�T:�F��Sh�sy�n�-5��&��~BRY&f{����l�b�?=��IW��e!���Ƴ*����)Q����օ�O(~:`U\��d����MrJ}"d{e(x�F�n�ڸK�o{Ob����$^5~l	��k��.�0I��.��!� �G 3nT���=p�����8�H�5x��]��|��$� �f�6�"� �X�%�*z�H�0H0[�≕k�x���;A���/��q�B�����1�����^%�ی�B�{��T}���ĞH��t�=��\��OĘ�@_�� ���e�� ������
r�`'��{�2���f��2Ty]�#=$�ޔ~u�?��8��E��U����M�ˆ���rl<E ��Kx�hQ��c)D4�҇�X�Q0@T��i�6�ncV�8���K�����H��Ut�L4�.����9�l�1�9&l�K_�<T�\	U.��<�w�����QZ=!��x�K��z���h�=�p��������G"�z��R�Q����`�ґe�Hoަ XQQ8�8w_rh�b%@�k6�E�v�E�w)1�i��e�w�W��\7l�ܯ��]�ᩆ�&��h'�WE�RZ��~1�Xצ���*�$��κV�?���?t����)L���%1�N�� �&Y�&�h��_\"q��F3B��K]	ؿ�3����	R�k�I� �k6�R,RY�q�r=����>D���
�H/�~e��}����o���(lv��D<�J�v��! ��: +�HH{�R;̈�|��#�gޥT�E�����?��Б+��E�f�P+;�����Y�U�M��w�]vU���MJjqeI����ޕ��~KQ�j!V}~��m�E8+[����%��7�M�6�!����Q"�Am�q��Ծ�;R&+B��f����$EQ�`���.TjQ��!ՙa,�?Ob��`:K��)d��h�/�E�㠣=N�S�00u{Q37kv1$��x_^�+��j.��~b�u®`���+Zoj6dVqE^h�9�x��$p�%s����њ�D��ٹ�D?Vd��]&b'K����&�y�(�;ܡ��I���P&
��:����^��D��՗i�Ĵ�k��{��������5Do�Z�Hmv$���v=�d*�Y�9�A��y����%l�\�q�٘4;����x"��Zu���^d[^��0�K ^*��@6���ܴ�}�Z����+�?Xxd���J)�E^ ��H�P|m=�"nᛁ'J+��ذMi���e+;���7��@�
�$��?_zH�Gd����,���O��s���V�ķ�
����w��O��G���B_�a�"� G��`��^KS�������-��t�LV#h)�1zv>�ٽ�����C%tX*�kc�bWMgf�۹�� �|��&~��I3�D�����E*� �[4�~H+�����1r{�l0Egdƹ���1�SP�UO�$��=��~F��o�w��_}7Q�ݦ^��������>�/��*' �_q!���G<7M�B ��qx9i��X�s��|��5�����ws�߲Ӗ��,	f�l�ލ�E:J�-�bj8�0��{|���Rs��`fW���=��u�w(O?��%,�Շ������#��K����])����$�f[;T#�Ǽ9�A�)"l�^�3w�W,-?F{ *��2s7��[ɼ�����I[���8��L#]9����i;+�4n�ʹ����0���)n����D�_�x�<?8tj���y�G#��b��oǂ��=Q!G�Y;T�QY=�_��Z��Am+�a��E��	vu>�R	�)=���=�49.99i_�PqD��Pc���+P.P�����AwI��� �/��U@��U��>��>c��!qW��%6���
s~d�K�������lp	�^��!o��3z�*�;�6���}� �=֦58-у%,�I�Ұ�b9��:���X��$�q�o`����nTwsGR��te])p�xj�	�!�qV�{igLb«��ufMw�2�e�^��>u��3�}<�ka��ͻr��XT�������.�Դ��^.r1���b�lв߻[�}�����Z��37��c�ΰ��$�+T��"+��F�PV��,�i�g)?ʙ6���a�̭%Y�z�k~��_/��~a[�R옖J?bQ�GLD��d��GlLk���r{�-S��U�g��K��_�2��b�ܒ�z��^DV���_x�	��N�$�I���󢡛�2�l�6M�^"��Ix=���}E��Ŀr�#��yد����	�����1B���]y�2zL�B]���f�S�3Ξ?����p��zs8�\�Nkzv]�/���X��8�؋hx;����c��w�<OS0F��������8(�T�o��{����EDʃ�> �6�)�`X�&J;%e���SA����d��Ăi #��Ϣ��7��%�)���vb��fz��/q@!`� B���� ��� ޑ�̬2K}�v�.�*Uڙ�i�)n���J��ҌXE�}�8R�IaŲ�=��I���Fb�3�� Hx���)���>-��4 ��3�|�ԭ��)YgD��{5t3�ŞՂ�����	��	���&!��.a������c�V�ߙ��h$pq@�YX7	G�|舖@*O����@���,7���ܘ�DI�M������x<߯�8.��f�����a����d�̟f� XXuWфV�G��Y98� ��	9��5����(56�t�վA*twY��C�"g�*�Y&=G
#��Js�+	)K�ƢW�wH!�8���1�Fw^Í����Vj:�KO��q�z�j�l�-�������0����*	�ŵr
��{t�eV�_�&��{b�tf�����Ā�"�דM���]�8�N����H*!�g�G����>y|����q*�@�QC�4�#β�o�~M���!��0�N�ƍ ��b>~Y.��jh�N(��V��%I� ���S:�z5l�q&�e�Q�M3~���ݨ��t�(��_?$��n�)v�~�v