XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K����F)Oeh�F��&YPN�y�o=.b$v�q~��^E
R���_.ڴe�mX۷����< T�T���`��aUl<�sǁE�:0�wfį"[�����NJ��,�E�o� w���l�0���.�xF�F����/�ñZ�J��q�/-����@~FF8׺��>��&c�޵�M�S�i�F�:y��'W,ۙ�<t
<a�ޣ(�G�>����ޔ-���]��)�����5>�>��_��#r)���c1ve�Sx�-�t!�ضW�����O��9�t*�M�|d�4QgY��͛bJ)��}x��/��fh�L�l���`6o�յ0����t(�W�y��H���>)z���r�k�B)[{#������>��5f������D[��� ǖB��mީN�l���u��>{z�6�8زIh'�����h��~﮸E��OK�n�q�6�-��H���3��3���;�g�����oW�&��Â�SJ�ޖ%�y�IQC��x�_��G�;؍�!j}�
�$X�3?t0o�>�}N�y3u�Wo�Oـ�:`rC��?S	��b���>N�A��Tz@�N� � 4� vUU�]W��v�u�}s�Y�� �j~q6"��S�闾4M��ՉD�A���'��v�t�@L�`=s�MH2:���F]����~y-F-3N�UF���P����N�e��ܛ�<�P�_t \hBcv��V.<�h���+�4l����]MG1�d�E#� Ÿ��x(�]a1��(�4XlxVHYEB    2326     980J�~��C�kP��I�?P�i�U��}&#V1#AJ<X��K�u~��(g��"��бG"�S����B�?d�#,��J��������d���z�q��2[z�[e��2�������g�����xН�G��r>��kV���Oɓ5�o�g�2�A�Ӑv��J���|�C�N�+2����@�'��Y�BZf��1��^u�A���DZ������`S�x#��jKfZAu���SÚlR4Q�֗��m8���'Z���e ��[�Cx�]�lbYp�P�,p��e��gV=��Yc����l� ��@��+^M�/B,������4��%��[�X���5O*4+�z�>�ާ}�4)�Z�� �C�db6�5_�K|�v��[J�z���M�{�A�p ��.��ŀk�}drJ�x,�0�y�YF��,�����ت���� uZ~v�"zq���/����C�� �Z)�ˋ�Dl�͓�(���J2v���k3����㻁��H�A�.�HV�I'��plH8_qC���E�KDs��ij5�ϊ�]Ӻ��,_��d$��R�+<�Z�f�z���bbJ�[���R����Ħܟ����LG���h0o:Dy1eY�RS}$�yw����N��u�}+�'%W�p�rk�c#����V����wtx��	�U0�J{�)��OT-�6S�̓����D8��s����h��Ҡ�����5�!��3��X4��|^�r0�����й�����2��#T�N��􉎥Z�Ojgsa�Bm��GzԄ�����d_��m6�
�1R�L�%x�HC����*I���c��e��T9��Y��fӢ9l� �>:�!/ ��G�/L?k�*K��{_�p�?�9�'#s�I�I���9|c�����7U"�����APơw�j��<�wp7P�R���v��������GJ���+��9�W���s6|p�ՃϚ�RV����ZV7�#�񜯸�?Z%���^Su��{��2H��@׌p�^ᢙ>��alS�]f���/3�L�'!�@�ˆ K���4��y�m����<�n�cG�[7PtHr�]%��+g��r^��Q">����h�|t��TK��!YsX1���J���Ƽod��9�Ŏ��6��5s��!i[�\�m�F4g�[�����={ {��B��.k�S��J�p�l���eJ��2@���bq]h߼`=o��<J�c"]ߍ
R�w���~tE�`�;~�d�g�-����\h��Ig3B��A?�[dǘ�sx�{�������[�n%����:���}<�����ܜC���c�- �PKX�Αí���B��Q�y���Ӥz�S+ӊQ��b�hrqQ�mg����gw��k&c��Y��j�a�0�F��P�������b��-j����%�V�E��L�3lQ�ϥ?�^���!�o���,�
�$?�z�� z-��Hj�^F�w�g������F`�	��(�6�RG����ݦ7�ߗ+�Z.༤�ڈ�D\�=賖9]ڷ��4�y0��rm��z���Ǩ|P��@DE#A2�;%��-�y����F��;^zX�( ھ�-S$XܠU�"���[��R|�[}�wf��g�������u���ӑ�}c�^�V��9Dd.��F�iȉ4<C�
�r~�4�*dm|�ՙ���+Q]L��GǏ�.���l��B��h��1%���V��7�L�C*o��r�f�����=*6)���Tm��Qx���*5�@�~�8�}k��>�Ħ���~q�_ٟ������H�<3�/�ƚ���)���> �7����Y����n��m_4'4�Sl7�o2Y^/�?W1���I��YD,T��Ѽ�U��G<�?5&�#��q՝�΄�3\������d�Z v�

�,V-���W�a�º�8�j���� ���+r�kH�������x�y���i���׸0�~�B��#�.td� �;�2���غ6`��k��Wn2�v��{h��D5_=N�����p����*<fHL5�_'4c��][:0���i�?v|�B,�S�/�d�`�??����U����r4�'0����r1����.{׀KJO�4��H5h���I��P�e�M�k~j�?n����y_�8�0P[�G|�Cnv[�\9oI�(��ܪ��v$C����p�� ����&e��A�#
��QH߰� ���(���(m�F�0��6�@���nH�:�T�]�⣮�r<�&���N�6Wͤ���tzƅ��	��&�Ε���z����p�@��n|q�)��i�-G�}j[�6P���VVٛE��D����������� ~ ��G��u|<��c��{�rO�юe�����|�Kd��5���Zh������X�ʐ��~n�De�3v�b