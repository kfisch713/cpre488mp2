XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dEXj�Eí�ጂ=�N��d��b|/�R�bGg��<P�ӄ7�t�c�%6���xQr]}9;0dҺk����*��)#rzt����<U�
�c��c�ӕ
��=1���pg�\��0�mF6�Z��P���: ȥ@,�@�it��:Zϛ\����B�bMs+g�=u\��'s�uR�C�Y�m���<�m�����-�@��7�s�؎�����d��?⻀/��"�]<>Jq�s��C��:�����z���{֐�=�Ҏ�A���쏒��w_>��x����h�8��H� ���b|Ëoi2Wl41�%�}$�Y���"���4��~�b�{�Nd��`r� E4N��,@q��c�Af���ͳg�(ȫI��	p����5�E�����w�w��{��T�!�=j�Onʾ>�Cm��*P�)TE���t�E")d����.ҡ�	������{@�W՟��M��nqi��ϵ��l�h#�a�ǜ0
	��'�k|a��Z�٬$MZ,#�&(����3+IE�+��Q�J�[N�7埉ANB�> �����?�"v�][Ƹc��'��u�"�Mg&Б�	�U��b��"K��F���`@u^��nv�mߴJ���j����ŧ�2�:�bA_ 䰒B��D�{!s��Ö�=WB��qW�ō�5~Mu\�Дd?"It�O��}�+>M��݂�����˾࿣����[�V^���qN�tKR��o~����g_}����T6�'Lj&hX�>:ϿdY'-�� V���XlxVHYEB    2b39     b10��
�'�e�朁��|H�b=ZE&b d~,�s� ���@�"��l'R��H(z���ݤ1���BH6�Uվ�4RB��c�@>OJ%	GK�5���2��L⑜S�x*�~�����P'3�%R#�e9="I�� ��8@�`��ܮб�<[�3�r�`S�� Pj�	?�f[%���BN�k�\�ʾؒ�h�kg���}W�ѵ��H�jg~s��6�x�u�R'=Yo�i��lT�G�	��tN?����~MO~8�x�4�N%���&�� iNZ����!]x���x�Ǔ����`U�q�1��qVNj-�d���{A>�	Ȅ�����R[5Bn"�t�V�H�nw/��8R&�OOQ��B�a$�(|��n˧�9��7;�E��\�i;z.u5JѰ��-�r��D�/��S�t���0NU���_��EiQU����i���S~4D{��\C-�+�B�qH���b��!�.k�f�؆֑�}N��rI�P�j������K�&�?D�v�'��4�+�7���d�T�s6]8[S�
[��~��G��ӵ�Bc׶�X��EbWg2�v'.����P�S=<a?&������rM9I�!r{����c�Q{��IBP��R�
�����խ� ���=-&V��mj�ŕw��,9w��2�->����� ^�X�����M�h��X���2-��m��*�0��\:�4 �m��_璢�Q�^��:��f�	�Y�I��c<6�S�_�?�Y�}Wd�O*�O��.O�\CҰ��Y���x�Ji�r@��y"�D����#�N�y�]��A�Mw;`� F�X^X�EP�ze[�S&��u�4�V������t��d1v@��5;����e;By��˲_I��a��D�͋�?�N�Ԣ�{�a��
2ه�{��T� �D�{��j%�gAo�m�l�����C�6	�D評
�Ί��8%>]�9�d9���8.H�̂�x�P2�� ����o	��!�̫�I�,Z@4n 	�N�����~�	��v�qG�vX������q	3�I3�+��D����vD��Y+&�z�YT3y�q�XЖ�0Q����a( �Sk�V_ɞ�����g������&��x��v�-��� ;)�ﰹ0P�Ƚږ�r���$;C~8L.P��J��
����������5��c2�E���Y�+�A��]�3M�9�1nap��°��g���ʫgƴ�E��*0(�uq����(����d��Iu_��G��F���Jw۽��i������K��u)���P[0J�.�Un�t"\,,�9H�_���I�Rjh�y��*�v[c��d?}u�
�`-���*p���_hH����@X��8:e\g���S�:��Y��|��Ӟ�>�1s7G._�q��Iw&��XyH��U<h�#�fUm0�JD�-l�x�Y�_4_	�~��8�� � 㖇��bn�<m
��K$��;HAj2*���xT'x�ьw� L���Ů4l��Q�Ϯ�E4�Ig��L=��F�Yxu;hlw��,��qN�	>fϳ1�B�<���3���0�+H@����4fN�-��V��&!�S�n^�a�΀������!2g����9_x�y �v=
K�/&%�&���:O�wZ� ���k�<[�z�L/bea���\��8;9�a��Y�U�2�@��Ş���An9В������B|�½�g`9��v���󒄅Q��T	b�l|EM��o�V�!�@�÷�E߳�DU��y�:�&�p5��M"�?��gQڧ�����Aa9zD�6��������u6��4�:.!�,+
C�6���X���-����oİw������u���u�t%
0o�䞘45�J���;{���QY�ʡ���YbQ�}T���!!���:��f݇U��K�⠡�ϗ^����A�c������Y�<�pC h���Q��6��XW�tMW(���ч�͵��$����D�9�)*��BZk�^J�w J��uO�b괆� �@�c`4�W��ڼ�n�͆����Tb��W`�7< 6��!��j�
��w����3��9���j�4��WD2�hWvfPx �t��i�,���H�Չ�ٷ���tv��Z+�a�
5�"�C���U�V�k⴬f/��o�V��6rk�b��l�߻��Wm`J��}�ѿ���OY��h bc(R��0��s�x�V`7@y�>�3�Z��` ^�ċ>�Y����L��W@=U?@��^�9�B�8��4�]USzr���a�.�C���=�d�Wo�M�5�_|V��9�Y>��I�U�G��Ů��%G�;�n�DO=�g�s�u�^�'fA*��v��hm�xR�r� �u�u�"�+���� �3�����gy�|�1�������g�Q��5G�T������1+8��ѤA�^��|�f@<&�������kd�W��+��_^O�f�#֟�rw5sq��%;�	��X_���2Ƶr���4��A&Z�B	C�?���VD�A
m��7�PYf��"������x�c<�cl��Ȁ���X��ۺ�x$|m���*a��gT�FVx%�/x��\�<���]��!�53`%A���Co�G&v��ST��>E�Fd8Zmi�m��'���h��_5�t4�C�v��M�dN��j�N���Α,�;m���3"g����k�N���n(z����c���Vl/AO�ް�hJ���<���������S^�rQ�_�n��Ee��b�!&���b���d%�=�)�Cj�O�\���cj�