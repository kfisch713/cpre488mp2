XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��؇�n���H�h9P��tQ3覉p�y��ᡰ:��I�6э[��7ʆ��ńw�/h�S;���1U��Oq����8�n�q�l�F���Vj�o@%jw���������ʼ^�P<���;V���С���~��R���vj�0�0���;�Z��;�`�s�ʤ}y0��) l�1�A�Y�y�_%�]���lX�B�,�֡��F�.?$��3���J���Gq���R.3F�Gգ�`�_{�٘�(�rmLD_�WH�i|��,kS���#}�X)�7��p8��Ʒ�?_�ԥ!|��� �6_�����,l̂��b��hbA&9��h���d�f����[���R�7���g�W��_4���5�UQZ�̅���U����;6|��{�p�� ����td��ӄk�J��#�m����'ɫR@�4H��G%����$����}���*i�3 4�P� KQSJ�����:�r��+�*)���3�6�W{�C����tR;o�V)��x�Yz����@�j髳��Go��nٓ��������ct{tX[��)YG_�a;��G�첱�z%n��5N���+&��"%�b����U9ox�&?�n���5�i�O[�9�J��.�s�%`V��lܽ�v�~�<���~�z
�gQX们�~��S�݊���=�G_	�mp���:H3�-���C�����2�,!>� �l���f�ԣ�`i2W�������ك������8�tc�[0z�8�֞[��XlxVHYEB    5224    1740��+s&��
��M_���nt�q(�pe�of�!����M�w1W�"����$��0hBN���!�n+�R~� y��
���DX���;�'�<����sF�|���l�!0m�6>�_ª<�D��g�6�Ӱ����c��gXW��S�ؗ-���Y���ҟ�(�$���ޘ�b9�1taK�����5e���/�4���v9��=�c�_6%�JslWX���3����Yc�"QW[�|Ƨ˨��-O?^[���b�V��6���ۇ�Wt��Z�����V�o�ه������3���I����S�tFQ���J\'H�����E-��5�˻�@��U-��(U��f��FG^l0���^0��x@��[�
n��7A���^�Z���Ǽ0��Q�;O�ҁ6�T ,!�b�cK)���F�?� ��}�&��j˝p@넣�,����fU��gRu�.�Į�wz�}�~m)?�&Md�lۦm��6F��v	H�������=DRFwo�r���-���bܠ3wVn���*k����'q큪��o�ɤD�x�*���^k��ؐ�ltMm"���<���bS�**��usH�+}(RAe�SH��/eo���0�܄ғ���h����-�|k��>���Np�o8��Ϙ1�r� ���y$X���T�:�az�4��&�e������+T?4�`h�D�v��#H������B��M����n�B�QՑ�y~ν����zN�&ή���������k��u=%ћ0L[9b$��QMmW�1ܲg��d�3B�T
�CӵQg �u�DN�g��R��c�o'�ʷ�n'ǎ��l�
�����eUT
̜0�T
&���`���P��P<���v�a�:�{,F7���^JD�WEL�4�k����0>!�i�|
�I._D_�-P��x(!�ͯ�i_��I&�d�����X^�!��#�'�V��pO|K�P�wOٖ ���$x�t�#�������Llw+Fdd}G�Ei��8��n��z���W����fk�זY�5YpL��uI!
�2�R��R�7Yx�
;T�1+0����/��# ����بY�����*�;�'���J������R��mH�N��>��yAO�;ґ<
Z�i�!�^&1V�}�8y�:{K��6���Q<Oډ�,;4Fӥ�_��6f/��P��:5�b\[�⮋��W�s��e�+�X�������;cvm!)�:�jT,=�Cˈ���L��Ю�"��5Vb��SA
�	��%zY�����EQ��]`�1~�Ҩ!B��Y���:u�k@д����;�dٿ�>��NO_����({HmrZT�7� ;F��t���%N����|� �H4g"�R�I��BQ�x���U �I��4� �s�a�N��m�9��d������75���y/�<2������2�xq�Q��z��5���go��nc�L;{#��eWm�H�X�,�k�#�`��["l_��,5R 7!9d) �v�;���o��!���Ob�q���@Xǚ Xg21D/.�\�k�
譫Q}��l�Z�[ ~�g����)b�p�22V�]��勏`_��������켼B��0����5���Q%p3U�t�@��xl��P�Lf^�!������}�\̞�����x�eI����S��������5��4a:�3���F6�:���Z�5�e�㖳�K������$O�:��KiHl�`�4˾���)i>}c8m��<��V���?̕ny�w�c�����,e��]���R�ѲG�H j=�&�#����rY�ݍ9aF�%�����99��6���[����Y�׹����;�k��*���,�=������ixi����֚�=��Π���(N��?!�GH��i�c���ok{�`?���W*ي��כ~I;lva�4$+�ID)�҈sBj���t|nj���<T���Aq�!��:�j��^,�]	G��2U˅���+Y�
�h��^��nἆ��{���Z���8h�|�e��Q��I9�a$�<�n8M�Xe�F3�&I��(�G�4jyƐ�	5 ��96�b�L��T���e}��ZU<Y����ù� �A�)l4:�N��<ݱ�o�eb6��Ӣߥ3�9�z��Tk:Q&X�ZA}}��?��{<7���ῌ�0��GT�3��n���x�g:.�w�{��%M^?bO/����4��Ӣ.�o"X�-2<GrO��{WAn�u���ux��[d��<I�M���6r�@�r2]��i�)������,.��7�O95�8�J7�j��]h@$J����u;}�ӥ��7�+c�� вL�f+��<]�y;����St�id#��"y��i��/���+�^z�0ߵ�-]HC�yg��ױG�u逡����!.�zC�e�8D�<�W�15�� yXj��9�\W�����E��i6_�hۻ�����߃�L�Ěp�8���u5��Q]��,IT8҆f��f�0`�aʢ]d�A\�׆�F�R˩�gRhNz��xJF=��0|[�Ѭ��h�jJ�Ym�I��A��xo[N*eh �`��8_"�?J	����s����U͛+M:�BƸ���SJuBLPR1R #%�(�[)�GT>U5���/a�l�YbD�Ty=�(;q���i+�Ȅ��
����Þë*G�36��JyX�^���dr}�j��TG
�Y'@M�3�>ȗ��s�w�mRY���u�I?j�P�X^�P;��*�9^��n&�>���s_K��RV|��^�ځ��-��(g�
Xl�Cl��?9c>oKR�\���8����ĝw>npݗ;���zNA���v\	��@O��EM\$��_~��ެ��	1��ow�k'�jE��;n �B9�]���kR��ݕ��ރݤ�24���@O�.��Lfbm�[R�*��)�������J�?T��bM�q^�0�x����5qΆHD��%����7"��X�t0E6����ȝȎ�HJ��Nb��[ͮFDz39-��u�vb�LV8Iٌ��G�y�٭���_Z�ϭ��F�^�b����4�%��VTh�\��U}H
áB�#}���ҵ���`�沅&�u��dtb������<�+��&=�k� ��Y`��@�Y�R�5�pK��~_�;>Q���=��έ�O+�W^R�k-v칧
����ܜ��^�H��N�f�����V>�_�_V!]�q�_�Q�C�<��ة�D�(�Lޜ�țW ͧ��(��m'�riv�ZY���|,Į5�?q����MPR >�POL&`�cuS�q,m(��<,��ҚO2��o$�:�rEH��ڻ/�6,Iu����<���'��@�"�"5����{Ao����S���U7HOյε�����������,�ߙ~����PZ.k�r�����j]|ơ%;�TurHȃ��IS�q(��Y/�	ZE��O�x�Պ>	D�J�)�|��}~��K�`3=� &�ˎY�l{3|f�����O9�_��)e$��HK��Q�u��uGK�6f̧�?����ce$b�t�\��
�` d]��d���C��=�����zk�����f��i���[,�F8A�Yj�c�}w��%%ڿ��+�Z����z��
}��M�9jr\�i��P�x�e�� +H�}��ݞ�\�=:��bn�(����j����ol��A��7�ЧV3�U��o[5�������c��t���[a�y��'�h@�� �õ�K�$��i,�]X�C�Hb�+MRw�<p��$�]�͸�w��f-M���L�tv9(Fy7=U%w"T���G��vB�e��n��+��Z�)k��ȏj���b*'V^G�P���ձ�O�qO�feQq�Od@�|_��<S�Q�!��'�`��ߋ�	��6\���=�{X%zte���V�TŶi��W���J����+0kg�C�����?�hF����W&�!�V�;����@�����p�H�Y�Xq�n�A��Tm�ҿƽ'��"�H����jp=�v��c	�>C���n� ��8ť%p�M�q�����Ղ��-m&�?+�sB,�:��_�r�9�0����Y��'��%1Q_�M�8�����g�+E0��z4@�H�vu1-��n����*����٘��
t{��6Ҵ���n��+-�@��x�ͼ,>��5�"��4�w��{?�+ ���J�5Ϗ�@��O6��b��²��Ŭ$8�4�Bc:��ط�_���u�m=�3��EQ���ƧM/7mn�)BA晵������;���-��}���a"�i�� f���-"�6�Τ���+�DC���
�%f�
�"��s��&�����F��D�R5%.���@�'?�`�jĶ�|OBg2WKS��I������!��T�����%F,�O�,*p���q�bʍ�
�.V��m�_`(�u�����C�����a&*[`;���J?�
�����_)b�|&F��sL��:r+��e��|\��z�}:#�x���]������4H(�%�����ѱ��|�,f+Q�����%�t2Z�g�K�\�/�v|�h�QdF��
 q��!m���9��|?0X�9S�	ZV��G�B�6����q&I�X-ؘ��,b1�x܄3d����4�W(R�'K��w�'��uL�P(h1��@�Il���Q�U�d� �(�^9Z£�_S�`��~��c�	~��G/�<g%2�/]��D�dZy�Jd��b������{��<�����}�ja_�K{X��C@�.��˻�MHo��!Ybf@|-7���qx�FS�Q8�K��Tˈ�Yt ����(P:���\�AEs���k�*Ev1U�>��b�����>f12-b���r+W=<틲v��r��p�s�?�>�6�==�Y>6�~۵k�@���|F�nX���g�0XN�6c�V�<�ÿ�}��=U�/u�_��������_�����}�:Bm����G���M<��$�7C��:#�f#�
Nh�\Du��.�s}8J�������{<m�ݧ(�4_� ���9���9sǁY��qhlܝ�2��0�t�!*ș�N�C2f8%ݯ��.�����<�ݐ����oٷLͥE���^ȃ����As�?�z�/�$��Wi�U���ˋQ�Q��w���P���Gh��`&�����x��y�#�Əyr�s@v�[9GE���VM��q�Ì}��$ �+q_W¢I�fSq���)�Y-c�8�Zg �9-�>Lذ��;.���sˠ0�	�j��Ԁ.dMn���j֘�)�,I�X��؆���R�ΐq��HK4	�^Α}�D��;wO���n!;�T�x�'4.�_�Ϗ�cV�0Qd��<4�gc��F��W"9�X����2+|��;#�S��H��Z�b85���f?P�r5F�	�1�j�b
p+bq?7�I|�JBZ,��fctx��t�灢������Wnt��=��$��'W$�c03בI��fY7"��I�J�i1#�����:�KWxc=^ψߣ!L"G�zD�BĞ��U��<�ˊ���r��^�bo�3uo�L�	�Q���S`f�������S��p|�.ǧ�G��x	�����0���u�b�)�y�ɂ�M)��V0��db(�T��l�����M~m����2��S~˨�����s'��g �	{nU�ׄar����Er<g��q��~>4�=�[3`q5�N�;q�s#��T����Wۈ0|��V~¼��Cu��Y�5�S�eY<�_>,�
�x�vIyk�[BЬ#�� '�mUęg�om��KP��B�m׾�� �fQ�)� ���8���h��ulkT�L�GX�D����\�yV��#������\�^.`�LI�D�R߬