XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�҅��,K���{�������M�O:%�.�@��`��M]9$�ݕ�R�͠S��9e���\���%e����V��Fo[�U�r�9�*���\:˦!���Fo�-t� d�?+����ht��|�{�s��e��I���, '��F�6��7:u5_! �b8�푀�F,�ꆀ��ݳ���%�ϑ2A6Ǘ�ҕ�8T
B��w�z"���9V���m�eN;3����֟��J�&H�����TQz@�;G�A��J� M+#`O\���wo�]}�5NS<�����B�6u4$�����x���,�AI�nf��x8\E=psV�����	�"c3�g[Z��n�~��5���5����5omZi�a��T���T�<��%��	P�	g{}p�P&5�0Y~/x[B#��!����!/����ҹ�c� %G�R�H��K�~�[�#�_�� ���)&r�g1��f;e�%�]bI�{�f[����%�!��k˃7�s>��R����7�K��B���(����؊�:x�Uv3�s������}��"�dx7ʚ��~P�h��r��!3af�r����YPJ9�������*�Y��Hg��k%�5H!P9	�'-���vaE2�9�l�/햧󓮂X����X�r.��t�Ȉ-�s�\&���	�d�72NтB�1���Rk�V!��@�	����z������l��c���]b�Ga���#�N�����%}���P��f�`6`��N����i��XlxVHYEB    4284    1110���:�Gt��4d��S���R3̓I���_�:�_w�H!�����]�s;*���g��H7V*&ʹz
�#� �<�<dw�`k?�'Q�&*�<̋�]�g[oD�:>�
8hu���*Bgj{6��C/�y��i�\����Z;�'��v�Os�7���<�d
��=����������*��/Z\�E�tS��m,D�I4�JIL-���Js6��4����Q�nAw79#9_7��R�\B��C�~�i�i������h9��(}5�l3{���S'ş֚~����w<V���[]V߭xT�Ś��z�,��)��w�:�3�#�ߔ|<��hZ���4�2�tXk����N��}��6��^Y1��rU�e�=.�c<gs�?m���$o�Ξ�A�������H�����9�b��x���k:��LۑN���]�Y�����b2f�������� t�3M�a�;[���C��y)��{X�����Ho�D\����ڙR�����}��j��YH�п�!����c�
��l�k��aA\<�ڍ :��� 6�/k-�<�h�"�%\[ی��?�px�d>�Z�䭁wPր���*����D��H/̡'ݒ������e��eP�gF�h��U�����F~��q��!���NV#�(e��E���8��2��{�Ҳ�|.L�k�;R��@�C
�r y!X1d�����P��9H�JD�渭3��r\흪q�1�������kn*v�	U)�<�/Z� W�|3��j�]z�c����u����wb+��F���,��t��6΁����.��Qwu�����)"�r���s@��^�-�{�����g�Z���C��(m:X;WbKrU��V�Y�0!t��ܜ��u(D�EQʉ��	vN,	�gU���k%VB$���W�:m��G�B�8��]��KP�,]yg�:���e��$�z �p���f<v��&� ���l�����~t���E�̈́����~}#y�aѭ8yѱ!H��������مJ��o����6�p��22f�e,��M�cA㲟� ��C�wҌr����jNj[\?)A��Ҧ��=U7Q�i�my�|h$���e'I�.��hT��:�%!���W��,x�}[T��:&@����d�����t�Q^R����<;_!	�I^(��:u��eU�<>��2h���B܂��nB5SeO����7O�+�܉��:b7���-2!�V���{��<���~�Kn��o}J��-q��r,��{ �{�o�N��f(!a�y�.�֦����.�z�Yn�W��] �(���EW�����Na�|�ο��i`��jS�T����l;����Ҏޗw�t� Tn��=)m ��Y����Cd��&�Z����b�<C��짩�E��o�EJG3�;H/����ބ��kk��q��)�?�鶒� ��B%��)B��]Z}�FPi�#d�k����ӱ��n0�7ʑQ�n�-7����-���Gۥ�x��mCF���\0q̳��O]��-֐z�����<��Q��� �K�{Y��8\Ʌ������=��e���ӱ�¶JKu
G~�@`ʿ�z�"> 8�U����
|���Fc��^�8TNwJ�������t��v*Fi�7g
�X�GY7e��V��]h��h�ߎ�^ᅊA
c��5��׬!�o�����a�;�El�����媻w,ӴqM�e�?��Ɩ>���M�#i����*n�?��\$��b� � p,kv��YS�@����A� (���TW/��q��E =d����>*����#{`�QD]���B��6�G�)��{{����~�$zqA��b	��n�-��?w:]�@;��4<�5��si���s�m�������{$�"<$�21
��l]3+������LAŋO5(\*��*�U�� i����| ��A2]�
�
�1�]�+���,D�*%�D<���7S�*��e	I��X��?}(�:���ˍ�
ZQV	b]A�8��#7`m��x�,\V�K�y�}�ݦ�@����5u�yk=���\������ƌ����=ށo���� A�*�cm�f"�=c�����B���AQ�65��*tи73JZ���U'��n9-��_������i�[X�Cn���N�O H�<���:���}`)�T��Y��6�F?��Z�/���*�.5�Uw<\G�u����1e�~M߶Hַb'�}����������I��:pK��]�%�#��b�g��q(N<�}{ب~�~n|����ڬ�$ˡ�<�y�
���Be8��kj3�+�)�pWb/� .�}��R�!�iu�
�;r�3Te��MAY)h�}@J���b�CI����X���)7'[�����HQ!.���E�����=|�����6K@�8z��
��f ���T��x��^G���1cT��lz}���<�.2 �X�٦>�T�[8��ڱ�b%�y>hٵ�F�5>θ��9�P����|����n@c�,�$��I[�%��?޴)�[�ӣe@@�t�F���#:*=�5vgyᡂ������o����$�r�c��@Y<h5��DR�0�gh��w��x%�enT
�+����ց��� ~�o�74r� qL(�%9�e�}浜��Ewu�ϴk�MsYO��=*h�|\od7�=O��Fxy��� �C������&��뗂Qx�	��i��F9��B()Y"�+�kL�]
h�k��z�-������CK2#������.��΢Rࡷ��e��ȜTչ|��Il�ɱA��6�H�%�>Uͥa��*�a�Aa���P@$!������1��.�~�������'.&H�����U�tl�i;���2�]]�+Z��+>�	��_�~��YlD1�냾S3��r�[�N�"Jr�ɛ{MqT��H�#�>�:�}Dn#@4��i���/g��5�<{�A���}�+"$��Zϐ��<�ͮ<4����m��{���Oy�<}j��H�jG��Y��z�'̿Z����МƧ-��04�%�Ъ�-�f%S��G=�p�#�S�	������	uv�P�U�>F�l���e�vټ�<`vlC��==�(,lރKD����M�db�� @�W{��)���?��"3<lۧۢw-��G���<%�t��D���xZr#ivX&��\�	C�R�l�g �S7��C��4�Ȝ�t�d"���:ۀ :4�:��Nv5��id��`��8����ƞPZ���o@嵍�4ml��|�I���Z��h���qY��L�¼9��	WJ������v�B�f-���NUK�Ɋlj���l��oc�56O�Y��x�k���;���hs�Ň4r���j8�\w��~㮚�����q�c\��:��XB܆�~�Y��k����cA�X%@�l���7��25�a����)���l
&V�fqO@\����ԕiʜ�ԣ�Y���J��[��0�Z)��K	�<v�KI���Z��8����U�Ss�(C�p8n�0��&�O�]�~mS��3_q�|�Bp��8>O��+��5�ZK���P-���O�]	7�'���y��Ӕ���Q�8���ᅃS�d��J��PC�B,#�����9V+qa��?%�;�%*�n�fYĐ;M��nd�)3;N�ゔk�N�v�Ş�����pl�n�Q�x݁ڿ�x�Z'����wh������k�52�-�>��H>��G��L�B��[}���q>l�/D�-���a:�GHD�'*������U��:B�9���M�y2�P�e��|q�a���r"�H�|�6�����xDU�r��O,���n����	�M�J[�6MnR$w��3������e� ʉ���3��w�
i�x�WB� ��̤9�$㷨-��ay�ۄ�.��	���Rox����+�sG!O˜�zL|�q���}.�٦�vG�
�]���	�'l���������S ô�"����B2r�r�>�=��n�� s���"w�ֱ���?�vϕ����=�_��y�c���Y�'�ĭ��A��A+/�]�W/a�ǩR��ҥZx����8D�A���t�`���=W8��P��<���8�X/EB\;7+#���ct���C�y�[�_5c�Vx��K�Z��
1�!f�OH��$Q	�����T?��n56@�U��"�H0}m�z-	��L�i-�Mո.� ˟�ym�o��0���b�X͉o{�<K��|�x��di�B��0aĲ�oՎ<�@׀���5#���N��(g�V?),�Qð启���� �\�Q