XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f��bPr�2�k�ڷV��$���bz��^�I�R�5�^Uu���>���},��y�^e㩏 <f�Ĵlܮ����S�c
R)�.��v��e�ό)� �ϸ{��EXҩ 穀mR"W�AO��"'=�QD�I�6���r��-Ə?�R�XnrAԬhLt�]n=v%z���=O(>���-�5�w�юMK̬�H���Ne fC��&"�>��J
���!���h*�t3��E�L]aj���D�|���v�r��Q2Ⱥ��z��/�R���8n�8^E]��[��n�C�e��*��l�ǁl'��?9��{�:yZ�G;��S�TF��1�<�[�h \.9�c�{t���;�#e��k��A��):��>3��`���14�âur1��,}s�T�Դq}�]-t��/���(f�1K�����2A����Q��Ν��o���S6���z�|�U՜��(t@����G�[�4@W���)?� ="�٪�p
��7�-��ƚ�*��̅���o�å���B5t��`E�/ɒ��1S��@�Sh4��}�,��*w��`J�h�1��%�z5�V��?�%�׭DڐZ�I�X��06h������5�W�{�&G&���t��$1���I�{��t���pd�Y���@����Rl�9go��03]#'X�|��-z��?� ���h���6@��mթ�7�>�P'Q���̏�a�!��X������9�_�2�ӯ��+�d�po(���d�Im+XlxVHYEB    5d29    1390���J�)X"�xwk��u`!��(;"=;���l��]q�㻋�',wò7 2-����c��}��8�6��������@�̝�#�>8s"E4�h�[=� TU	.�,w�����|�,��ŒN���~a���p#t�8{!2���F$�>$ɚ�j�΄(�d�H�uLL�\X/�_^2�T��,o��=��B7RP��)Ev3v���ew��.ӌt=����p*�6�@aP#+�cJhq���xq7�]A�Ir��k �h��M�Y����@��I�-���"d��z�d��[��QЬ������y�� D���u?k�ױS�����ӑ�<�Y���U_�`7�*R��ǈhY���@���������|�o9|�h��{o�(�%1C5Q¼E�y�? 9}�?ʭ^~M�� ���q$s�^u�e���@��h3��*�p�:�_'	�7շZ4�E3�7���,7PQJ�[`��R��ú7aU��n�~��Lp��\�s��e��0��v��y����fM��JA�t�A�(
t��K�P���UfM�<r�y��}�&BH'�gL^~�b� F��#~
�+c�!��	f`&�[F��Bl�2������Y�78��~�H|1m�v����zBzt�;q�ճmW���P�+^�~Z�R�^�.��o����i;m�~��мZ$��#ɨMnC${P5#�e���������DkN6?���:�ݷ����:��Ȉ#���I8��jI�.�H��D�N�5�p��W˯�b�q=8cnbu�G��h�To�l����>T���5�U�e]Β��e�j�m��8�_�+����6�'4b���JÆ��To%�{bu�� ���.r�����y皣��q��T���4�/*�:�˘C�^�}"�y¡�U��u��[Ԙ%����b������G��2��~�2;)4Hg�Jez�J���  #4A�ȏ��>#�o���>������L:��l��-ց��P�� ^ט����oV�ǯY`�[��;IX�kiKрv�q���6�n+�+C���Ϭ�	�Ex�NIW3>MFg�c%����:�T�Y��Vʆ5b�Yr8���?V�g�Y��ߨ�)2���y�Y
u0PL}��$�F���7��3�Td;I�Ϡ��ntSbJgN�Ux��X����r��*Lp�)cIú�C�K�|Q����iI�6����/��q��0oJ[dlwgl��8(��ҙ���`{���q!��?l� Q����U��S�;�L�#\ބ�&�Ͼ���\�0F<W}Æebm�`,�>C�3FVZˉ�6{�߃�l��P`q�}SPԤ���$��0,7(:4=>Ux y@��S��b��<;��I:�L@
�kQk���"b�>�+�ʿ💉��A)S)ɺ����i�b�=D�p�;�	@��T��I�J����Ir(��_��C�;V����;h%w�t�0���\�#����
bIt��u��(\B��|<y�N��0�A׍��x۶M��~��%Z����u��[$� ���H ��2���~����9�Ȑb�z��V�?�Xq�9�s\��&� �xm!�B
t�`cHo��G~����'Nԁ�F�_҇DF=s���u0�u�9����:F�gA�`.�#�[���Dh4Vу�Ck���dY���"U���*С\L��b�o=L��U�����Y�S��)nu>���y +��Z�0�;�y��V|�9��Ǳ%s�7 b�32˼2	֏C[׭�T�	���H���7|܄�uJ����d���>F�T�I��nܧ����r�d��h9������:����[�(�\]^�=�j��/�,S�ǻ��D-�!j�cn)����X7��(gki_ܳ7ͬ���o��z<{��S �ݧY�%BM��~/�<?������5�?�/K�0!p��Y~4/��5	�&N�:��G�n��c�Ӿ�R�1�qsL��AE:{����?���	n�C����H��J�M�D>
�=S��,>q�Ro�V���T�8us�FS�[�j�+1|]+���(èW�c���P`��:s_�<��2p�3)���5B���-�-��� ��+:q��]
O���{�Q�u�L��ǴA���3C�*E�S�9�XйH+}�;~��z�ä�e�}?��/����5'�l	 [�#�,$v��\9���	�� �x�&)O���V�V�g�Y����Y21Wnj4��$���Ƣ�����w�%ߘ0��>j7
��Ä��:\!�h\�N�^n-o�@�W��)d\�~���6����L��
���	�)?;�~V�M�\dkY� >��%%�;����FԩS��0y�A ����Ƶ��+^�Bz���IS�w���"��;�I�T�Z��dG�DI�!�\���M��Ӫf��1t�1������ko)A ԗ㾜o��qB=tJhKpPG?>z��?���w�@hJ�P|Q?���D/�T�ܱoq��Eհ��sM`5e�L��:�=D�*��5xģ�`i�{f��kB�˾�؄ V�ns����=KN̥��}�Zhq��8��jG�v��a�7ѕnP����@����k9BǄ��s�����`�B	D6O;��ފ�E�g�ܜ�aS�!�\�����<�����d _��ʹhe
y�?�=;�7�c�(�_�푇�S<��`���F��2.o88N�]#@��35��ڨ^K��#�3X��c"K���`+J2�U>��Y���^:�L3�b1%Pyy7��j�%"<����ץ���g�o��3#m�g������^�e{�[�p�*�^�V�O�0<Z-#��U���۞�IǱ��T]M��C��}l��>>��`���k��,��u��@[8�D����z�7N���U8u�k��h]^����+%���J�w?/��4jj�
Rkk�O`�3(�ی!�@����!VʆҠ����^*Iw�$0���� �p�ʹU�mϺ�T��Ң	���E�����I�w�4W��1E�60!�	ei\��
���3��:�&��*��SI@��hE��O�f��^9n���.H���vWp����%�L܀ՍX����ě!��R�|%Z0*�%y��D�mВR��q�5y�@�����.��_V*�"��M0�g-S�����b0mR\o�@�]�5WOo�������Lg՛�W�w�X�_�������$��(�x�����ض����4� �J����fţ�`�[��3+3��H�9+�+��78-�P�3��21�g.�� *L�c�@��7Rb LOkr�}�T��K��W�H_��]�JY�y2��d�[d�ī�NZ$#w�nZ)��בl>����j�~1��ş=���1b�Z?(�A�Up[x�@6~~u'��S� %KJh�[<ᑄ�^�xS�^�:o��_P���<m�k���MN���b�B,�N*˱l2���)�;BP\�e�@\�)������`AIO߿�j�5$@�bI��}��@�R�y���W���?{�B\I�Q��z�na�@<�0����Ú�"�Ǥ����胥��_�Ҧu��4�*�h|Ga��Xa( 6��w��96O-5��l���loHU[\m��/�V��W˳Q�C�#�a"��F�Q�,��ы ī��o-w)ͥ�j�ܧ�(����(��+$�+���Ep���,�\����2߹dTaX�P�¶���⤫g�|uW��:r�&y�&��B{݁}�;�+�;d@3k���X��+��R#="R� �gKA�iwR�ɷoPc#s�R�G�V}�ڸX�����aRҍ&ʭ�+_o�O%q�N��z��3��yFZӅ���:"}��V����³�����7&������ܼ6���q�_�LBy8yq�l����h�̔棉! 2̈́_�[�+��
�6Jd��ym^~�%徃��N�}�M7�GiV��!Ȯ$N�����D��P)�'��}��2�yYd%��ʓi�J*r�L�z:��A5�����
�+m}�������ګ��_XL"V~e%ل��͜�r�D�$˿s�����q�u�]''���� �du�U�j�,r��=v�?�}{;V��0h]�U���@�H�7��'J�w�痢��4�}d�aL&�>/�@�h#h��l��^�9�h#Η��B*;nG�T�D?���[e�|+?"KY������5]�>�(,�b�q�0�}V��=�\g��y{�zL��-o���k�H$dq�nd"��&2礟w�2͔�����"��?�梼�� Ń�(o��\��)p�U�cz3#G�� 'V��*'W5VEⰏ��[
p1�a���L��<��ɔ���U�!�[t&���˵-�!��|(0~ia���������V��bk�h(�ö�Z�r�=�<*5s�Ӧ�ĵ$�_RF,��-���~M_��Mu��e*��Vn�ڶݎ	����Gc�d�m����Ӑ�-�_�n�Lc����-B�[���Y��G�p)��o�#$�����-Y���}F������~��m���`��N �Q��?�czJ��BK��:=e�]w+�)��x��{�*i���_ h-[�˽5s����}���f=^�e[Q�u�&ݯ�O�&Y����e�3h�\i1�"�f�������������`�<�}N���5t�Ť�;����,�_2��eb�,3�t0���x�G@Ȝ x�1a�ea��D�G��Q�7bS&�O��j�jyWݤXr����/ ��Gq�E��͜�����ȧ�B|ZABI�p��h>�崕���:F6�h���~�!��cWʢ���QM!��P���������3֊�U�����d�4yD�g��vS�Og�������EP�O���S����S*���DKۿjG_� dSh*"�R�晎&�un5��`9i7�-� ��_�A�]*�+4A{&ُT??cy�m�