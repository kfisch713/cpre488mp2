XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��tK-�-�E+�-��B�+��x���c����}�է�1� �U�.���F����r���a�+Y�H�)�1!�nk��Z[�J���%{/�����x^��U4�Sڌ��@����=H:5�.Б��O�QZ ���̨��ܘ&>��v}?Q櫾���ѭ&�TDNQ^���jWX�;�ĩ�f)Š4���b)L�	�,�w����B$-��H��
��rb�T�T��I\.�U��f����T3Rͨ4����"j ��^W�2��a��/�3��J�K�}����5[�
K��r1j|��Y&�l�ɸ*�ˎ�P�<?8.f�n�I����-��5G=e]þ���^��L� 9�l�ROg��l�菉����u��Kd�}�ߥk\d�Xi�V���y!��l��u�KKM�0���Ƶ�-mW���Q��	Oǁ�"�L>�c�Rrj�� �*�S��O�/ܬ.�&n���̥�)����ǻ^RQ�]�ߐq�����pF�Ymc&�Fb�FwB�k�čy��6-�1����&�^���󬱟���]��n�f(�|���s��{�$�żXH�#)fq�s.A�.�����J��p"4���7
s�V`@��Fz�O�`�8��� ��D"�hq<�����C���G����U��&�𾈛��[]|�|���ȲC匣 M�i�+L��@���!@_/9�x�Ύ*Yô�3�K9Ͻ��wz�M)��-��oo��`c�H�U��XlxVHYEB    6315    1790I�P~�����Z|)�F���:�F��0�C鈪�,�D�U�������g�>s\<���CEJB߭�ז�7f��IƸK5����6X��'�7���.?����"��ط"��Pt9	�oD֧��`=nԚ.�-�P]I���>l��p�uH���9�٢D���sg*��Yq3�Fy�`�	l��"Ŭ~ן-�v�@�(�Z��.z;SREq�xH_�Z{dU�` &�d��݉���C�)��Z�s�|���,med@����r��8E�nuP6���'9��CD�sD�w%
��"ti�R�Cw<G�]ݘ�{��˯|����3m`�!Y E4��O�6g�[kw�f��!�֙��T�W~ y$d�ڬ��4g��4	��P��sq�t�7nqy��G���Ψ6�n�-d��*|{5����KB���WaS;�<��m�?��G�����]�ok����M|��p~��y�>�����B�1�ǙbZ`R]6�F��nQ4�GJ������+0���R���9sXv�u]��Jħ#eHj��9�����`���XN}[E�[Wf����*\��T�6�j4t�u3�� G�QC����ܚ� )YL>2�A6�9��7�XU�lG�:[������|}�R�*�aEג)��M�U��>ې��M�w�1�O�=,�dѴl����=������ղ[����A��L��b9,Ip�����D����i*��q�q)n NR>*�xs�n"U0/���������޸_IE�|z~�G�p_�m��M]�Z,��E�F��c���p_�$��x��@l�\�e$ĹЃ��^���r ]
F�?w�}@Ի��yh�:PM��v�/��	��F�߷������H��\�sx���Á0�S��8ۅWׂ��&h�/4�P�M�V&/�e̙4ͷ��u�C���n�C~���*�@����V������6�����1�+�l��	H�.w��1Tns�/2�U������f�9M��H>��; BȮp����Wd��	(�/s�x{�G�59�X;���F��/�l7�z�I�>�Χ��wK��-ۥ��>\� ��=+[9w�$���
��[`C:HQܦ�L��@���jV3�{�P��H���Z��W���3���Mq�s,^{?�s�I��-����s\ث�"d\����n���9��¤�'~�૱uϘ��)���0��>'Y	'^"}�uwg���e]n�>REп�����4�j��D*!be\��|�.�+�b+��̹��^�ɤzU>|����o�ac�2_��³ʳ�}��հ%3?���dN��3����2a>��?{�.�.�L ו�
�5��UZ�xpt�Xh�CU�j�C��^´�?{Q7�Y�eT�����~]7�[},�Ч����L�װ�ԝ�U2�5�hA`�#�^��F�s`z��� B�q\&Y�6���#�P~����K��R�L�m�iow>���o���z���]����� �V%��A�єV����U^�J����B����WVNquv����bK֣(!��P8��t�Nص3�(����m��9=J��h�=GNVÙZ��錌��'gY���T*��c0���[w��������|��Ƣn.��@��-tJ�1����}ٌT[�
�VW�A��
X�D����z��+�E��F����`u�
~T��B�����t�n�;mL��� � J�� ߋw��:��E�SiG|=)�cU�y?x���a��0v]����b7C"�쏵�Ĕ��8PA$��e!�.) 嗦�,b+o�\RvkK=��X?�%�6F����,�y�����d�y��&�oy� L-2\�0�o��������R d{?��$�O`+�jC�hF��=�c�	�.[�$�k]������F�_�A��'�ѼH�ϕ.�V��炑��u��M�}���>�:,�li��^L,H�᜗뵨���+�޶/w*9�		,�9��#8 ;�|�i���Jn���#���@E�4�Dӡ�|�Y�sb��:p�\5��p�q���	QK ��+j�44�3,mh�FFx�k�����>�k0�9P�c���|�E�2��PR�eZ��s1�2�~�(��X�k�+�q�#0�:�򵀳�R��6��>d�b�Os���)U5�'{�]b����%��fi�&DȌW��2�'� �cV' ,s��
x����\�F�����xB0Wˉ�C��ux�<[�L�K��G|"�h���D�fa�#�\.m��#\��)�k�1 Z�,-�[��(�����T���a�6�����~D&�p{�2.��:�k�q�=XH�w{�jI��pG쏯6�*�1g�A�~L����������)����t�`/גI��I��qAT�Ҙ���>��,L�_#9>��ܐ���B��Ps��p��,D���H(>���G��_f�u���9c0�T=Y��1����b6f�Py[.��x���#~
zJ����c�u�R���]� :�/B���sخ���OE�)��N��D"���L�y�w��o9���;<�k�#|����Z�YH /�h$��u�w1A��	\�L���6k���� {5d$d|�ڞ>K�/S}7%OW?�4��a,3�	�ɷ�%�������\Yp�wVe��g'��[H��T����9�<jg��8�1�vAC{�/;�$f&H���/�2�t�|��X�yW(��MØ��@��Km&m��0 9z�Tl�C$��7~�I2��Uf���@���k�Y��
�Wm�L�*�� �S�����mB�?v�cװo{�y3��¿7��O$�B�\�"�Lz��ܠ6�l.�6m`5�j�j�!��1uM�9�1�&s�Z�Z�\O�(�n�tpG8�k	y�1����dcp�,�k�GH�E����=���_�� �#��r���r|i(?�+Q��D3��w7^{��9�P
�N $�}B�'��"��U� ���&"����1���EQƜ�O�Gش�.�����=���O�}M��@�� 9��I�ţ�d廹�چ[��q
ы��ew٢Y$x��������7�m�\�_���\��#�41NLXd�x�=����\A�\�!�M�Y�e����[L=�ƒQ��Ojr�Q�N�V���Rf5�Xj���bJ��+��Ġ;5�������A o��7�&rqQ��֠4h�:����e�8�I]zl�����P���;I��x�Mh�*l���x�W|Frj;�h8\��Bzi����#ԫ���<���y�d?� Hq��+�[_a)G�	��\aA=E"V���pT��9(aR�R]'/��*9�>�-;��<�H�\�3Mc�ּ�1>�mKO�˴i`����<H�����PqOe.��$��`��׈��w�qew�nL9�yг��ϰ�(�zwxڱ	���:�/��&�C�=R�pH��%*>��"�u*�ƤU���^���(�F<~k�o�����o�
ʟ���	� ����,�ܹ�����)T ӱ:�J[+?�=s7�h���3p[t�h���n�q���pN{�/�,��MR�$
_��b���% �9�4Ob��l�ń ���4edF;_&�_���1���Gd��E.��z��G��D$���:��W0�C�eM!�Y�9�V=9Y@��%]8����(�N�<o�s�!P ���8�;���"`M���?��w��f�����Ckni�Jq�8�}��_b&ZW��-�yP[^�����KX�#�m8����GXT?_��#g��-�A���o�uI�x%��L\6�]��y�l�!��N�F�5=���'�pB�0����Ҁ�2;G(f�)��
J\�R ����i�AI��\�!(φ���t>qyB�d�\;�E�$��E;{B�!����|��=���J�ț@�Z<(c\��Z:�_�E��{+�uD�*�2,'ȵ]lɎ޼��3�"�$�3���؉?�o v�/�wpD�
b�0���c�cK�(�[~�hX�52�/�n��t�I�P��K�H��������4(�����ٽ�˽�*�07�p}���ԙo![��U+s��x�l�����!����R��t�L"8Dφ3�eG�Q"(i��LP
�l��%��d�G�����	Ӎ߾Y�B��C��3��&�MQ0�uˡ)����b㺲d��M��4t8�x���X; Ʉ��*��Վ�
�7�n��4u � Y�֘�ތKI @c��Ҵ�ݱ��Jh��Ȅ�� �1�03�W��ľ�ŕV�)8��K�$6VFuZ����A꫇
�	`y�Of� n\@)0���d��u	�"f�(77[N��ɢ ��~7B��e[6�=7�X�
�S������-Q�����I3s��Vi�g�s��(�����$&���<Sc
��������ν�{H�'�B�Ձ�n{i��-�1��4�ұđ���GN�l���:�L�Rwٞ���l�63f�i���v�S���й6$�Ś�G&b���(��:C��D���� m'�'N%�)0��=AP��}%<c�]1��hۂ{����WbM�'��	ʾ�C��w���@R-82�b��d���Ê�����޻�>G�נ:�IG�t!f�(� �2�γTY���}48O=wR�;���N���� ��6�B�k��!z\�(����;�9���u���0��4�-�rl<��~�9�!�L���ܲM������� Έڗ��g;�V�\:Sx�xQ��n.�o?y'��~3�*)�쓅ţy��Sp�3%�N�3?���q�%��ֶ��}��o�F�!�܈?��}!*�J�ü�gɟ0��zk���Ⱥ�I�2'+��չ�`���YL��a�}�%�L���3`��^�����;R������+�T��:���ET���/V���V�%�*s
�^x E)Ǉt�F�\�5:8��E�x-�}S-9��U�J�L�X^���kL��6�w�H~&���gg�n�1�V�ox��6=��վrMyD��?g�M�TY&/#�?�`�S�b ����\��������bC��(h�@L#4Ψ#P��`��&�?�A��(T���m�qD
{�pw<!W�"~��6����hH���G�L༔x|"�u��Mg>D���F�9�$��Y�<�����S��<.�6q��T��c3[�JC`�־b�2� ��:�1-]�r�R��P�Κ����^G��jĵ�}�t�Ok40�=ЈT�kd����U{*'��p�X��Y(�Jbr�<Sq�'lƚ��C16b�p���?��`����A����ɼ嘍ғ+�+��'��p����'Y*x�M� � ��0*����F���u�N��a�좯+����xK:�h��SM�������"VX��[�����v��儎�h�C�&y�z5�uB
�Nxٱ�Mp����h�<�S5��n�Y��nU����Dńr�%�����â� ��ȿw�)m�^CSVod��S��9)��|m��06ހ���gxoU!B2Yz�l�I�>0+g� �W�N��٬���Ξ�P�eGh�~{�q��82lL�T� �L��fiG�c:��
W���&զ�a��H̓����*��[�ӳi���n����z\Y;��y�F���^32�e�{ �<�1�M�JV�#�|ʓf���@>���ohl�A~���M9�����/����gb���t�7:�=��.Z��1��h�T�΄V*�f��K��(���twQɇGo�e�7���u\�x��Ă�2�[O��?G�Տ�m��4)��z^pм|�X"+���Z��+t�������֐�p�]��J1:gC��:A�3*���#F�2�3�)�9�`;�x�(�@J<id�@�����U���,_n$$Rf��Rscj^�l��H�h