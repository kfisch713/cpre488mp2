XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:O�����}�?9�QAEy��:�}�?�&�`�����3p��L�`�VE��%��18�z����"�����x}�!>�D7]��Ȩ�X������,��;��JUn9���m�СS'�DF����ϧ�3�Nl���&ԃf��`�����&9=����P�Gc Y�]����*F�Ă�t�A�Vd�FXH�0�N]	�骂����7�t��gՑ-����J��%�<CM4��{�ʀ�R��`j�ɻ���6�b�KM�19�L	hǐ8�>@��{=��g�RT��{S���ߓ���3�'�aR�%��������ƜO)$	�����"�3����;q��T4�cðO�0��t���}�f��f���sS����L57i�~�G)�f�t��`���u�:�]�$��I��P,�Ɗ��@ ���\��ͱ�f���,��T͹6|F��WŜ�_�����Q4g���5މ���u�~tJY���B�����V�� <,�ԮCϔq�I�����ķT�1�<lCF���،�^��<�g�V0p�z�b��ԥ��cָ%�ܵ_Q��C^@��>����"<��Y~�{0-�%��1���J�&qd�%Ǯ����F=���1��3����9�b�d��a��ݬ����rOh��$��>��S֢�B'�uh����ߥ���?i�Ay(n���;�M��s��(c�y�kH'��E�ZvuY2�2�֔�|Y=���T��x����ߜ�XlxVHYEB    1847     900"�N����b�{r%J*W���5�Yx�G�X�%�M2�e��s~s��w ���ɫ�K���T���R�V�|�X�`xӞ7��V�gaq�Q��-�o�a��i7�&D�9߂~�@�Ҙh�'Z�v�+a��N	U\�'PJ�suq��
5�-��K��D!G)3��~H���tƵ���2��$y>'��"�ږ>3 �3�ϸ4�Z� ��3
�Ql�aJ��\ECV<�BQ@6|�$�縈����Kϟ�CM�?��AsB9�5Yu'�L���^[?-�B�p{D.�[3�DL�K�+;e�Z������7!*�p��[.�7T��MTp�6?E��g;��/;������۵q�^O��Fa�5o���N����m���V�N������~4�r�Z(�О=��Bm��4F�G]b�~aq��T�dw`��fGj��6�j?��Qo��Gˋ:*[�rk5��;�|��r_	�>	�v?Lut�	�ҩ����T�H5_����d8; �sw�P��}����}�B;tW\�@���/������vȎ���g��o����A6�����=��)�'��"�Rh�	�7��i�\�z�Fr�ƿyO�3I����������=l�P����>�F����be��N����:�m�TlC���Y��!�Z�.���h��j���j	�(�]�W"�"����o��Ao
�Y�XVw�d�t�U�㆛~���_0�DU`ӼG�@����q���x�d����ʆ�������mÖw7���?��cI�S�5�5���* D��0�J�z�tO����$D���b�����"Ws��G��)g�y�-�Q(
�s�"��>l4��@��z ����x^��N����S�7k.������N��8��5�������Y�T���n����΍���\��q!l0�	����K%�m��/���dGj�v�L~y�ֆ]��6]�lMgn}���,`�X��������Z����|{�؟i���k��½��ZΆ�<m}�- _�'��������b����~J�/=�x׷��ޜ� �?�(�V=�?�˯�V7d8�)P�r�>��� ���O�1�\������(����[��e��3�Aw��%�2��l��|����)�Ir6z�C�J�u3��[[��~C���@��^���3�e�#>��$}�O>o"(���2��n���q.��k��k�Q�i�{Y��	[��)t͈Rof4�x�w}X�r��T#5���atTY�[�2��$w��PDV"
\��V�Jh�q�֖���$�m
�X~�gp�3�M238�WP�nV�8�vc�,�F�G�W|��[�Y�J�>�⟄�-�leڒ�7����ӡY�{ŧ �,7��PҌC%�!3��
�#�+$=�>`0�	�Ni2^�_�4��l�n�l8�D�;�O�+z;>�D�0\^t�L���?y4��״ ��y��	��k�%�<!p�k}C�Pv�.F.0��9|thb��zN�C��bE�H��FR�t^���S!� :s���mB�K�t;�j��7e#áaCO�O[��ȑ�
��e����E�^ʱQ^�F�\���z�'�c��������<��w"8(΍���d���F���A��X7�"��_��.�T#���
��s�8luܘ���Ճ]R":}�60m����oČ�N��ַi@/����c���;�0\���a��C��V����v�s?�3��8@w�
�".�:�ʳ�L����+�c�1�4�@��{a����T�cCH37��ly��g��y-In,�n��.+�hy}!��Ց!����R�Cr����J��̞�G;;B?"mq�[:2��~҅Xw����~v�CQ�!KG��t�u0]E��3*>(������W�. oj�f��J���b��[��6�x?�c((�f9^aG~��&����!h�6��w��Zˀ�+��\�3@^�O�԰z��K��|폠�C���m��}�g��ϯw=X��w߶Շ�و+��ڧ���o!T�����2�x� \���>Pcb����`�V+E�G ;�H	m1��Yl�M�Qh99 *Bg����n���2�f�
�g� �F�6)���QI����k�x��w��,;G�j��˨���AA��Q@��j�=T��c� Ə1��p�|f���9�1�g/V�M��k���v��z{2"!�e�:�OnTF��5��ɻ� ��1A��H�����y�p?M.sI��z�dq�нe!6���
CDТ�@P~Ul��