XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��߾|�a>�o0��߸]M�~���!k��:l9�ݙ���)g?v��2C#��#��NҦ>s0�]E�a���}�*��V��	/B�u��|�û
S���lH�r��Չ�ûT�k�X��dr0ɢ�w��S97�?}t:[*+鰲���J˱�?�+}x���\�{���	�1~)�!��U��̐қ�^$׆���$}��
&��\��9٢��qfm^�,/{u �Y����5�@L��+�����'E��Io�ӳ�i'=*=@��q�)������~���&ڡ����<��R�:F۔�H_�����M�V�J��Ad�G�A���|���7a��N[7���;�AQ9S�&_��c�57ƲC
,�F���?���0Nι�l1G���m��
��3�e���k�@P�����]!I��*�w�*�Z<	�h���Ѽ�s8�/�٣*~*0��?b5Ngs k
�wK�ֽ�
��[8�a �����$��k�i�$2��&�g.�F�A�|�۔�`��j+=3@��w�PHH#�o���Or� ����H��K�=2��·��dQ%]�hQz<�J1��d��a�Nv6�1[�I���������=�p��$�\d:��tb����� X�v%6�e��#�n$C�R9��XJ�9�����#o�ت�1�X�o�\2F������C[E6<�đY�]^5n�"�2����Ce<{�E������_�#'�7Pd����������
x���w�;2�z�uXlxVHYEB    5cad     f00� ���՟��R}-4;E���_�)�nqT]X7��ǜ�S�E	���B�\V��[L�%!�b3`���?�$$^����)��th���2%{���
�����ά�1]]�� �f��[ǲ_p"i!��XT��J���4:��\`�CH����Q��&�U؄�쉀��+U��Hh�m����ٵ
�=�Ŗ*�M�>�!�Ĵ`x�`f�=����ؼl���2nb�:�	�������w��qb�/�9T�����,��$��NP�b�X�c�8Z�$i�X����X\�@�wd�X�j?�q#z�\׶D�u��F�~�.�\~�t���5�&�y�K��y����Т�e�`yI�nb�:�G[�P��>�{|�G�T��}��HT.ǚŔ��=�#!�P�4t�{�g6���@Q*{.���g�q0"
�ap��Wغ.�_]���q���צ�XM	�� +8���H��+�c	���`�ǎ��XoR�/�BC MQ�o��i��(��9!	�}�Ѐ��!��Q�v��r�R����v1��ړU?l��oh���X?�ו��F	��K�I�ϑ����*�7��@�{�z	pGq1˪�ڀp :��h`Ic��D���*\���U��U�`jw��4ٲ��,�E���K^�ȥS����9M������P"��IT��1@�p���w��(__��k��2ƃLP�(��>+�����*Y���'��s�x��&�S�xP���o{ f���f�PGeg�?��E��|��/�{x����S�����J]v�1 �`� ��G.,�v&����eC�6`HL���;��X��i1��z���2�ja�w߶�<�Fe�
g�i�N��s�9�ځ%�co��cI���@�L�#Q��5(KQ���=of���o�Pő�p�}�1H��z4};�g��>��nШtW*5��9�~��3���gi >!�{�te��b�ۑX]�����4M0hT���X���Q!��0���#k]�p�g��$rmD�r(���U�FU����}�^.�"!s�]xiy�OLyO�Gd�{�N#��}� ���X���µ�r�P��BH1���L�v�U�Ѭ4���v��N>a�u\.�2N�#���v*t��%�.��9�W=@DRB�~�z�FEITw7�BKg�
[�Hm�$j�ib�tz����ɑJ�[��493��(� B��8�æ갪���>�N��+��QU[MO����%ci��L����WoÅU��6��M�S[Q��̟�J�i��*①%��?u�1��c�Te�~� r���iʕ�X�0��W�}:s��9��6��`��i0@�~�t�
���mX��*1�%�Ĩ�sb��ysr� K�ݏ�* �Ðf��~%�@ۅ�/����~��^�U���{��#N��8$��PӪ�����$54WA��؁ai���M�[��=��>�e6/n(���~C�t��z"1a��z�Z-jN	��:w8pk�x�nn���B���c������D׿�v�Z�I'�R�I
���\�����֒Of��vL�bT��d���e+�/�/'����N����h�\N��|%\'���~ˋF�m��,��m�f37"�8PG��F 0]�=J3��ZG����#dߞ�C�}�M��p@��  �Z)�B�󥘥�%J�m�oXr��a_�N>e�����r�J̚�j���aQ<���n�nk�
{2�Y��q�[�tB�g��(,�J*�>��a�辴L{'����X��?`�Ł���q�Ѥ�b\��TF\o5#�u��Wa�hjR=W®+��q<�Y�:������V��('AM�}u)}�ԁ��H[5l�P�2�&3�-A����Q�/.8k{����Y���="�Źg�)Vn�Ż6�D��[��Ig�*  #pY'7��������#���SK�p���!��.�8I1/�Ph���
&�2��'ڳ�������B����.�i|VlwX1�+�#�>q�'��JU����2#K���3���O�'*8u�V9��~M��*�� *��S���!���,ކ�y���@'�e�}=�q�_-٪o	 ��O�kZ�e����$,]܁���10�Iv7�l`�N �<���ܣO�>���m$.]c�?��y2�o�Xᱝ����Hb�]&*�L9��z=UX����G��Ԝw[;���7n	}WvѦ$�������=%�V ;5�6p�a�
��~�?�*�*�P�|��$y��P�Սf�o�am�VS���b�����m�a�*��5���%��W�&�uJ��M}���d��c�)y!����䪱��9Y#���E+��#��v�/A��a����T��D+�S�����c��5�讯�+n���%���^��f�d�+bQp Hx��@�H�/u�`]�&��a�x7�$�� ֭EX�	�h�K���U@����h_R��~XM�f�޲��<��b!Ȯ���������f��.j��ŃK�|�~ �rkb��%�?��2�?(m� �6(� 9�U���t��R�/+CKA	���ww�f��0�����t�*V-߂�\�	�S��L�J�.�E���>փez5�^mj}����:��F:}�=����1<
|s%w���SZy"F�lo�f�YwI|n�Q�7�Me,[�:%La���m�HH��8�ke�B0�1ܱ
���2=�o��B���<s��_;��A*�Ѵ^��;�p�8����L�7�(�YL�8>m��҄-m�{ɾ�PY@�[]�^N�$/�'w�r�g�t�IV4��\���
�;ApZ��D���D6��c*�n�Ϗ��b����Kg};q�Vɿm�3B��<1-�iv�gieN�l��'K�y�
k
9�ȩ�	��<����ıp�s���CM�UGr��(��j.�?n�z<�a�5~�KU�
�&��V�nS��ӡ�d���K���{6�����ʗ/�)�c��g�3YP!���Ѓ;�)��\3�ܛ 1���Y�����ɺ�
N���_��0�3;*���b��쒝��Qɢ�{��A���`�p�p��($N.���������cQ{��,u=@C����L�Q�O�"+j@�Xfl�ɇ27�O'�dN���7G���4������R�[�џ�HN���T�`�d;�C��*eJ����� I����gZ�ͺCm��H�JD��!�9�h�r�6�i�Q�֮��T�H� k��qut�E��g;*0��T�!ӻ��KԕE��%{7&���E�Wj,�kP�G��6��&BI�<b��'�2���B=���K���h��o5 ���Ƈ�l�[��3��� LI���#���C�����`���@�y�©U=�p���KGO��+3� �8Ŝ����x�Ѱ�c!�e�T���)��<���+�گ7 �%���xh~
�l��Az֒�Cl���:�hŨ28{m�^S�}}�V����K��*4�."$�H�DT`�`*pc(��6Ȝ��ok���eI.���p�8b���,d���1�?�'�3%�\����E�І7ݰV����Ӗ��e�y=AiaIV����nHA/s����w C�ί�9�A5�J�ˑr�~����;�7���z����ޥ�����|W+E��s�Tk��F)�q��cg��)^��χ��CKG#w��0�A�BJ����KTF�E�}�k,�S�U�D$#Y��]���+�ƺޯcQ\\�̄׭J�j�B�>	;Kc�m���ƘL�6�/��4��{����.����ȺUJ�