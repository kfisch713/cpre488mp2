XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D�q|�U���=�hk{t
��#OG׺NZ]�t�2N=/}^���C8��_��m΂�̉CV��oW������([��%�B�#(�%\�Re��&��q���0������n����.J@����R�[Q@��3/;���䝄�$pUX)ʢK֏.T��2C#���ת��n��RE4_���y�I�x��
���D�>N.
�a����B�b�ge�U�A̽\4��".TjnVO:B���b����Z���i�|�K�5�y�QK�����	(��)x�K.�}�M�)���$
�֔�u��-������������T��K^�ѻ��P#���.�D�xKd6�IT�)�����̧5I���q�}޵�툭����]�ʀX���C�w��h�0��|����z9>�yB�5�������F�)LhMCɨ�~����2����j�Ù�Յ�O����b\�L�%W��6�A
 ��{;�y�(:y�����Z��R@f_��]����st{����Ã�R���aAL�=Ey�\!��f�2E�;�,-_ya,� ���l��|"�X�V6E���u!g��m�*:.'am��ʂk��d����Ė�h�M�k�_lq��=B�ld��@�&���VU ������8������l_t"-6�x�J���nEP%��X����D �����FQ��I�E�{���vܜ��0��=_٨��F�*����؊)���o�g�Qe�;˘���:���t�XlxVHYEB    af58    1ac0�ޠ5�8fz��18�^-GO5)
��-��D<>� BбҦ�L��s؉vm��L�U2<�Ԕ�/�9�3� �
C��6�AJ2����=7vh���:�"~x��S��7�,���f4��7]�W�'����E��Xp���<?�o�RCg�W�y��# �� �M�&ϭ-*����poV;�˗>�G�?.����+�"k��Zu �W!�e)��r�0���Ol�B�x��g����������~Ǟ��e�O��ߟ�|�ޟ�R�f?�U%u���2ʂ���(.w���i�{����ǋ�[u:I��v��'�:4 Q��H����X���V3x �s��7J���!Q%v9�s�r�H@����~��e�T�=�@��l���Lo�ӿf�B;�+�����I:+�sFA���9�$",��쒬'���e�A�c���P�z�T���Sy��0L=�"pc���=w��+��hy���>s�	�r5���mI���?Ň�q��+�s�Ke{3L�T
(N��Ԩ��ҔHe��pݰ즕�]��e.	�#�IX(����4��<�\��n�}@9޹%������w��ͧKD]xxeɘX{ZS%Zﻁ�j0"��Um!�/��Oj��Sa~�^�O���s��S���r��Ze�O`���V�AE��~����9^CTW*�`rT�|�
j�4��l�
�l3��p�-�������/ħ�O�vl�;JSD\��5*-ǃ
���V��b�B��Y]��Ȝ�u{�-Nҿ�H
�'OK�}�����[����+	��8�:1,s�T�NDka'}}��Ǩ�r����ml<�\�Lˀ�&�߮�:�R�r����j��ʟW�ѢJ�/��Xz�*�2X�AUeܢz ��5�cC�x���i<�> n��N)�}b��yݲ�:1WA��8�c�(T��*��)�ۖŝ�!\9�ZA��Qm"�Qڏ����T�i�]��9��bb��8���ǳ&9F@������L�f���[���0ÜL�o��]�nXT��F��V�F\!� I�"�(����0�d�F���X��1�*�*Q%�NG��}'��x��ulEȬ�0rԄlg�WFN5�Gx"(�q ��N{Co2�K�t�Т��2�`��.;R^͠�i�����*Ѳ%xD���|�{
f�ׁwF�4ݳ�o������^;&��Nij`?��QĹ�ڌ�� d ��U� �\A�'���x�9ƌ�?Ӫ�E���nk)��X�a�����8Q][��fH��.�Z�VK��a��YX�����Oy|��*��J馊��25Yn�G0�_h^܂���)��k5C��s�r��Z%�5�&ؓa�=�RҦXu���(��"�j�V��Q�O�mDD��C����(���ov��r��=����=�Hߐ�ɖH�l���mA@S���(��d���K����4:�pi�%�tےO!u��B�i:~^�Tɼ&(N�[�(u��
�FO���[�/�ps�Ox=���e���*�{�G��E�=��.
�M��xd?��Ԟ���xy�H�L{��)�pe.��Y�"T��P�����_�ɪBA�S������\��+�\�5Yg6��Q�� ��a��>#�^ɼѫ�,�h�H t	!��s�.���hG�^m_���tm��=ӏ�d�+c~7���sJ%P��w(�?��a+�<��\P\%�	�~�@9g����a�]W�Ƃ��	�������ܜ���	�͊&�1�&���z)B} eDwiyv�������!m��fUs��l���yp�Y�M�\��Ɉ�G �V�Ifw۷��&o�"���Y򴃓;>�BC~QN�[�8-6ˆ,zt��j��v����$�5��/=.^V���+������@G-��!،Q�)33.��9>��3M����ޕdg7~���q��_tF�"<y��h�A���m�I��ǭc-4�a%�[#�[��Eyox� ����g�F��S=4����&�]LWdo��P�D����H�W��Nu�?�W�H��|ocj��q�a��a,%�8H>U����>��_��Iɺ�L�Hj�i��_&�Ѧr�e����#���4@����4F���ZNs7v�XeF�U��N��B�;��GU���O��PW$�u�\�Q�'Wc+��,25'�P��d����ד4��3�O~��h�:�:	�z��x�<�h��&�5��څMV�A�ʱY �F�3��)�̐�L&�>�"�M�qp��)�����P�ݔ?U�}��+Ʌ�UF>{�h�F��ǖ��b�n��\�.1[:?j�2���'v�� � 
�I����7�-� 4��^�;�Ɇ^�����+�W�n��8���Oi������ת�0OL�&C.r<5lo��,��j
�H�2vk/|��?j�+�۳�Yʤ�^�o���O�+����
�t��� H���z��٦9حAFU��n�Z��8gk�<�2�*1|�P1������ȝQ��,a�":�Y�w�&�f�:��6B���,$#�!jj�n1R����eX$��.�$��[�Fr���M��R���M��E���g����X�nY��N��)�]��0�C����0��VP���2^w���R����w�|}�ǹ�a�ڛڽ d'B���JA��F�z�x褧���F,8���m�q�D��C�� 	MY���_x�{b�����lQ�>T����~��ᢔ+��N�
s`X�q:��߫���� �b������]b����qyȄm]����3	F���3R �ڐ�(��29��6�5_��@SτG05O��<Aj�P��������j�G��n.��v��iwAє�XE`�n��v�j#����eW�W��,H�bv�P���J�z(Ŭj��ڈxJrj&�	�(��'Z�&C���m����	On5&4�����ޛoa��ޜ�{��� Є �#=K���q��)������$v8zZ2�
�m����d�R��f��	�±jC�G�\�U��T2���v0�t��f�����
y$H(���~]A�ߨ�D�p��Y\��G�@hP+�;�d^�z�47�i`�}~��w�I����vQ��"'�zoB�:u5N��1�X�KMCQ�����5r�.td���Q����:/��q|�C>�8�d~��au~�K-d"�y���@6�! �����?�]�2YLLv�p��Mx����������ƣ�RxǞ�u<�ț����v���;v������z�V����Ȋ�F$�5�@P�ĦU&Ě��a>��S��4�]���;|L��E�vV�p��&z��|@{3��q���Yy�i�m�:yz=-Õ�Y�����G�_�e�k�Պ�<�Q��yU�
O��f@�{"�L����GJW�ȓY��bڝ&����=�!'�.�8�sL@�F{٥����6@PjO<�[�r�+�V� Μ��������ĜmY�?�\�T�%��ƣ(��d�m�	/+����8���z0(��$κHK�.�*��@_s7�ݧ�v"�_|ܙ��jBf���i(Q,|��m�9�	����Y�T-�͝�
l}~%�;��=Q=�_�c.�l�Y������,���X��IC���T ��<4 ��Ӈ:�R��ݳ����*@�5�S�VkA?�sdR�pi�0���cӹN������/e�̓�.�qΥf���&3]�ս�X����q;2�`sq��{�ǧ�lX`�����L�];���E&���q(�9�\-��ywY��t�nQ��3h���(W�	�Zz��v V���6�eӉܒ��W����e���IB�<_���'Ky�0����'�'�&��0g�s< @��[��Wg�ڟ�R��ʜ�	���c�Y��V���� G���}�`��#��j��.�JO:ś����\US��+�7��{��k��2�n.�]j<����
�����������EՂ�S=5�1�5������(����.
��@��JO	N�w��y+P���Kˋ�9d��8o@��G&2)2�x�t�_�&�g�?�"D�T�h	<f2q��@�č���f8�M`L諸R�y1�}�Xغ�` �q*+tФ��u��)[l,��G2\�Y��	$e�KoP��˿�����m�\l/��u���ah6��F�^n�PN�>P�9���۪��u6���� n�$rZ~t=f�ƚ>����F������ƭ3G`�_�y��o�>f��5�:����-w���ER�q7��X#�z@:��k���0c��֫�5w/�"�]��o��߀�o5��������.���Iџ��8J�����:��kx��������*�F�ő{ĕ�x�G����W�oI}֤<�1�����_�l��F'
o���=9r*�pV�K�ZԼM��g��y�J"Bhu �G��T7q����;��V}Ӧ�䕖%�P!�"�Rd˃��^�(��R�@[_^���qr1T��X���	ң^�dbW�'V�Ț9�8-<�[b^���_�A@:��O��s���iht�\6�FT��*c&�%�����!�ִg/�}�֖��	`Lzu°��\?:�>�n�_O7��7�1��x\���.)�@[`��,�l�H�����r��x8<��1�19��R���f��Է&A���@	B�5�o�J���
��[�Zp��<���G7H��A�]S�}�Y��� ZF��Vזt~4���P%�E�Hᢔ�k��ý��mA$�O���%��/��o3cXC�Hғ��̅��g��ł�q��%[h3�z�j�_�?�!�-�6"f��X����V��k��0� �Ϸ�pdl��	�7k
��z�/6j'�ek���/2�͵#;�N����Wܫ�\�-X2���F�g0S4���k�>��&��n��f}�
�x�����0��TɅ�ci�!�g�)���b#�X�(�z�o�s�`�K�^����*҈��S�s���L��?��螱�#�E�y����8��g�J��kʰ�X�X�I�q�z�~��<$x� {���8 �����[�?���"����7�^�ޓf�͝4�.����A��"f�%ܼ�7��fZ9,�Ra��g�g�Nc�E�8{&O��L�X�^� ��&Zw�ӕ�$7�cbg4i�)L@8���e[O4�ƿN���7���|y�V��6�'�ࣈ���_OG� ��t�s%�4]1�޾����O�p"�U=]k��1�9��z�FPڼ����ϻ�ƒ�h�Q��8K$��C�0�;�#���%S�"���	?��:#\����&�x33��6�+�w�����|���V6�|t���;��q	��N��|�3��:	�T�J�O�Nz�ٵ����y��3�ҩy��q�8Sa}kj�p.���H�ǆ�#~t�8s�4L]0�bHE@ �긧PQvl�dh�]��#��_/p��kI4fL�3�ځ9=����I}�e�=�Ha��LL��8�^I�۳�6ŉ�5i̼����o���ۯ�p�lbvE��*��n��G3��գH�yy�^��P`�����'��b��5w�����`�l}�lX�y�b���5 b���_���[J،��u�:�����������0�����h��j���I\B�ҡ#�����{����T^��hES.؀e�]��ؕ�{ >�?��[@ϼ�BsD���4&�H�������(�۱0��d�	F'��fi$��K�5�Y0&��kcCJ���2�x��8'JR�v��ԭ�R�K켯�����Xl���K���M^E�܍D�@G=���+lv$��0o��b�]`��_�Zә|�3��k��?�_���
��$:���]k�Y���h���ߧA��J��1%��-��de�~:m��l�t����)Z��2�7��h#�X,��}}�5l�0�{�:׿ٳŔ��A�,r������d�b��Ľ���Fn�e�-6p�ƃ��lݎ9��Ie��������,x�r��{�]c�c=�h���L�����*��<|����M�|*@�U��n�`���.�k/�1��00��益����[<����_B�6�J��⹭��`����楸���5l�'�؛NQ�Lt�cm�v��G�'߅\��&�tsf((���U�O��+�.�����N��­y�E,���9��~��		\��b�Tg?2��+6M�i����ϝ�%Uu4�p���Z6�0p�^��.�v�>h�p7��\%}W�	�X�B�$
ô����i��/\eU燑>8��Ə���#YF�6����/��9(�j���CiWbO�؟Ĵ���
E�}�e���*�w���r�����RL��a?���/�6N+V�9�=�'��f�
�fj��S�'����?�Gd@q4�ֽ��z��d$S�W.hD<�$�6�$�ݣP3%�I��|&@e�zF�k:3W_xƴ����W{W�J���b!��SG8���c�WQ!�<��7}�U^ �듒3�f�B����n�K����}���M
�����7���~|g��T!!{�]�㢣�������b7���8��s��!>���d�
R_	����T��.��=Qx�Q��q��\���P����,M�q ������A�Qp��48��x��0���ē���q�6pʦ��$2�tpԧ0��`�o�3Q��D�<��񵶴,{C�fJδERc7�#�L�[t�a��k�(?5�}