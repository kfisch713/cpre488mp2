XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������,oӦ��ԇg�q�Um���ϕ���`�9��Uj��GI$2���f���S#�2��֊�]���<Q�`Q �Ľ��07��o7�`����C�n�D�>D��>�ʂ�'�0��l�����yo��.=D�Zx���a����4��9@$Q�,������sN���ȯ:���6��F�<Lz�ō[��#T��k������?PFZ�Nj���|T��=��i9�}�Go���<��9 T����8��KSxt
NV��!G�7W5��O���x�?�5�e5��oȝj��`���5_�w������mm��v<��
B��7~�b�1)�O��m��"(�E���޿�H��n!K�Yl
O�Ћ�T) `�|��U��GGTfE��f�sW�� 9�C�|+PQr��a	��<��v�r8v�+7yz��<f���G��N:lv��>����w��cU4��~R*�&������5��x���8��=�'����@}��#����SSFW&Ծ&]	�:(��h��{�[�-�R~n� zݶ���V����u>bQk��'�y_��hV�6��ɨ�2.���]ب���r����3��<`=��3G=U���g���iԏ~���%Z�b]�c�{'��U�v5t	�ł ���( ��8l�$��fXC�5xO� i��O��3o5����em�Bt�{i���p8Ѐ0���ʄ�Yz<��B�԰}>9^�$949o���[2
���-�XlxVHYEB    9fc7    1fd0n�b.������og^�ˡ -��K�͑4���˭�|_�ţy<蘛lh�1����Y^�]ݢ�j���YĴ C���\�o�+�W(�~�;���"�Ȥ�m
�֛�y;�,x���`��=O�R��|��v�Qq�pv�{���4_������(q�ԉk�D:�����a%���2�5�X�H��%�+��.Ӈ;��?��ɽ��N�՟�&��֑j��+�
B�.�<��¿��!��oB=��d�xek���$��eVP$i�X���	jN>̹�S�W}<q�._�4��{{K*X�+m.�,��`]�B���#�(���a�n>Ե��uE�<mw��Y0�[�W�R��Ѵ@ie����h��WV��J��4�UR�VĚ�OI�z��3률�PHx%��Yd�]����?I@+�̺��7�k��R�����;u���t���A>U#��s��:q��E
��7g��b9�%[A��P'Z����YU�����(��>�=I�}�]�F�/b\�)�h ��lj<!Md�˧C���G���}�7	Hj�$S��aU1�`��]�1[{��)Y�aLK�라�G��<ʬ=|���
}rk�m����U_����8ަ5v ���8�m��N�L/�s��2Vh#��"��Ƹ�/^~��/t���E�O>i=;��VjN
+%eȆ׺T1\�\$����W�򤇨��.�s�� ����S&o�-�@�ȃyܐֆ� �Y&���BW$̊�Y?i0��9�ڧ����η'��_ݶ9���nώ����������i�1J%��+��E���nO]�,�"���O�T�h�DCfm�����DCTz�J� 6]�7����ʂЮ�ڐ��愛�,nWY����f���iԩ�U�{OD�b�q�c�N��]���Io�Hʻ�I�8�Zq"��9k�WC�:��s�����I��РAѡ�1��ɿ�6Y��Y�!U�l���Rb+��$���{���\k&dG���e�;l�e�IF-{����䃖+�Jp����i��8��t����Cܾ�0�[��y=��N�������0����>V>��I�Eb0����U�\IԞ��
���.ί;��Q�r_�n�ܙ��N��G*S	>�&�Y-l���쨰PM���W�����mH����]��'2p7��&̪�=w��S�v���^�MA�Nʑ�T���G��8���%�o��2a{�C��z�5�ؘ�S|Q f�f�o���d��ewqG�s����%�16�}�x�s�9���LaD������e_�߷�b�Zh��C�G�nvD�p|"�3�J��jq �4G�#�RU#�e���×q׈��sw��wD�Ř� �$\���dw|��<���n�m���`�q��Z4�5������GF�5��l%�WK���$8G'���ā��M�%���{쑫$	����a��'�i��z�ܜii��� ��]A���>�{��O%'�1����S�����bm��W��ڱ�Di�K��& ���&MЎg���%�3ݾi�0~�`�'~?�a�[7^�B�0��H�n���u�!�Sė;kϐN�jP߭@��Q�d��5Ѵ��?릹��9�~�'�d��,kFʞ��IFq��7�JP�D����kѣ���f˯�؀�Y>8�q��C�=�����s��~5���?~�����d��Zu��� ۥ�aaqc�����i�Qvΰ0J��Ƣ�2�tJ���)�+��	��N�d���񑽷� ��goCz�`Q"i��?�$Hl/�Ҟ¸Lr�tm�o%?7���> �����]�()�c|�/�_s���b���e!7�ai��~�����EOy��+Z2��}/hR43��_ti�z����w7ȉ3a�?��N	X@oR��~�~_t�-��V,���Xlu��������v�%� ��X�x���mȑ#�������Rn~�i�D��*�>�J�B$�q��,�Ct`J����ڑ>ӥ�4}�����cT -�xX�c���X�.e���TRY�UA(��~��i�͆n��u�s!���q�awB���`�{@ω���l"+j�^g���D�qN���"X����E-b_�]Z����xig�G¿^IH�b\ex'���a��{1��D�����n�͏����T�f�U�Xp�tA���Eˡ��Í��-(�i�IW��&��1��杕���[C���l^N�T��
����G�D�����{)�dtG�R��u���//�r�BvG�;��8�����
����KGiC�H��d,�N���s���y����yg�9��H*v�O�z�K�.�d��'�9Q`W;��͊ut�˹V���)c*1��g}�@_��|�5�W���C0��� �5)1~%}M�e��S|����;�sאPU�,�%���H�ҩEۆQ�x��m�]A����ї�C��!�p*�^$���-�`5> ��u���{4�>9#X����R�J'b�W�.e���cͳTbЁF��u�M��>͡?�š�HF�Zu�j�>���
��4�ϕآ�s����A7�-߽x������צ��h�]2t熋�w+��X�a�gc��(e/߾�����~�Z�O�A�3@½�L��8t�\|yv7���D�D�?7�؁k٤�"��M�xw(p+�ֆ�&�戡`#ޫe=H��}F�w�1;��`G�s.�}IE������g��#���«�U%����Ѫ�a4���D��G�Y���m�ƙ"�> ҡt��j��0��e���E�.À�xp�-�����q]E���4b���,G%�n4�o�}���^��W��9[����N3�{����X�V�����/S$��S<�)�d*<�l�).�r�%����٧ÿ�"t5)���9���)k+a�w\̋nvάe�"�7�:�� \���a��-��9Zb��^����p>�aE(2HQ��7�_�x�MԖ�0m�&�L��d)m`��,y�����;���@�j*�|q&��Qa��ҙ&X��~���wD��_���F���>���V��eɯ]%(���>v�{l`ǟ�e1��<)r�,|�&�]���R���l2T6�w�O$��*�o��!u8p1�Lk),q�^(P3�,��x(�Y�k��S~[�)�s벋 ��1�q� 4CͰ�N��>z1�w����≃�F,���O�z���"ޗh@��&�{�V�fg�Q����A�TF��
�'�]��,�!U�%˰����A8���H&;���tv��(9�A�����t�ʐ|5�׹J�'�Uё�N���`܁'�b�Ͳ���}[��K�Ae�Q��]~A��:'��u�753j!{��b�;˄:ƽI���I�f(G�o0�+�Wi�w"�"�-�aqI�1���/6%d�/T٣�쁹P�� ��dR���?
Tx�UR=�Jo¼����Ŝ�C·��]n{5���C�52<ޑD�zj�9�xԽ'e9K͖���o�9�n��86�4�D.0SA����t'��^��A�8���ޝ�af�3�o蹽,��E�j%����Qx#?z�ج���`7G���nq6�
\�D�o�Mt.%-�lG7;RLlN9N��¿��pO�/Ĺ��R��]�V�xM�d(ʘ�sG��A5~�M��j���ꫲ�R��x�u�S���^Lv&�`����~����9����s��q���j��L���n�U3UHuX���y1I*=�\PGh�מ�������t`աVu��� 7vЉ��\}��	�0p�����M�!m�'Pg:�0���~-\2��]0�p�uȧm��:ϲ��i�����XxWP@����w�(v�/��L�6q,!�$p����g� ��?__��-��辀5�E�'f��b*�@����@O�#X�ժ�=�4�gٜ{�8�K;m���;����"Γ���tk"��0爏^�}�݀�J�opuԉ%&��^����'��9�:�0�9>��Hj}Y�Ro���ו�	�[�7�+�o�?"EΥ��!��E�3�ښ4D�C�pX'�8D�ɱ���oۈ��?��EG"i��D�'=�Ƴl�i�w�k��&X�^Q���t]��x�/9��x&c�f��Zb�[�F�A4k���6H��h���v���tBq�!)��M���+֢�?��}}���A�����L��B-
ř��������N/���V����;��s��G���<3�B%A\�8����y�[�t�M���i�S#�4��(�"%�3�P����Mĉ�0�o���Vo�5�����p�I��.�i[wym}�{��PEY�&_���:M�~	c��920�8�h؊����#ZƧF%��Y2Y�y�vX�`��e�w%���8ݭl?�u���47~��_v��8�+IB�q�@0� 
����N�27�����\ڮ����N���B_�.���xu��fڕ64iC��feeŝ�5<0&��w����ʑ�@�A�����m���n���j�[S��BK��U��v�s�x[����g����l�gxo��Q2s�7j+�eI#[-}�?{�Q��zn�a�u���ܢ矁vS�����ݸ����]mL�Svͫ�jd�馻��J �t����5���]��q�6�}�6�约qxc#�<��"���Ĵ!��cn�8z�����G�l!̿�B�"2/�U�$XZ�S��[�weY5H��H푵+�!�zhe45� _�rV�;�gQ���Q/�P�U���:v��F�aOu�_t�h��~t�N��.)�4[���q��*��E�Cx���hq�C��8��E�&�3	�.�)0���ֿ ���ҏ��������^[O��<��(x�/1�F��p�NA����4^r閧9o����2�I1r��)mq�S7��:.��f���O��uD^�э��~�J�K:_�K������6&��*0��YcZ�d�句Ai-r���_��Ք��It%jtQ����^F�I�l�kf3M�J���kh�N�%P���j�oF�nW�3�Q0��w"+fObl��L�nŵ�~��0�ΆMg+�����x��(�WH�Ǉv2\��)����8<�}���[�oK�-u�74��w�|\�0uU
2B ��&��b�����O�a�ղ5H��ʲ�#��_ �aW0����B.��n�3}��V�����mW4�j>b��"!߁��֒��aٯ�D~Ź�;��hʿ)�Vg�;D)����!κ4���cq��Ւ��*���B�w/�U>K%�0�^��)��Z�Y�Y�۠�d�p�{>�]�^J���U�=j���x�8 d��b�V}��)t�I�+�,-���.ׅ�ΔȰ]P�8�)��sQ����2�r��u�%�E�H}��֨Z�|������A���I�D*��S �rO�K�$�C����(|~��diH�_�;X�"�.�a7����e���{�� �u����O� D�2)LŻ�b��s6Y��f��*2�f1�Z�կ�+/����l�ʚ��Ӈ���c%_H���W�͉&��b�v1ڭK}Ejr,q3~p�d��~���Pޖ6yt�nw�{f5ʴ?_�}n��/����ߙ�^dRd*�D��+%\����t�*�ujv&eT��uMrE����%G뚸.���bڿ�L�!�G�:�p��}.��~�cbmyJJ�Y)��,2r�k�+J��,ڻo5��m�`����{����K�B� �L�sM|�;G)_��M�4��֔� 4r �X�������H�;�le�	��D#N�SX���N�KG[Lk��a,�Ż�����篝�+f���Ӧ\���`�0 �ѥ����6�\/j�\#���^ź�D�� �q�J?v֘���1���_�G%��E��I�[6�\�S;Y���*����5�8��.�9݌t����|�F|��R��Z.HNĻ���Ƞ��ŭ��G�UG��M� ��j�9�!マZ! �ݵ�+=]C�:����%���A���:��89%�����^���1���d8�G�ɣ��޻7wT����A��&��XF����������2��E_bŎT�D���Cl_6�H�Jb�C0�(�b��x���UD���d&"m['���~�l3����kTӼ5(9�'�:'�XÀ*�a sIpۓ�g��#pT-vS��б5��-�ƥ(\LbՑ���z̫Q��JN�_=}$g>�@0�M'��P�2Dj}���n�Pj�O�R���	����x`�>M�KM�����謤~����|lLA?QXq����V碑3B]c!��
6�.8�(���5�jxv�:`9A�P������-A���$��'z?׀g�ߣXB
�T{H$\���?��/�������l�9��a�:h5���΁SЌW2�'��cݸ\�C�3]ȫD��X��䪻l�'l��73�8��L�h��'�i�?���))b)S+�s*�o"1�����h��d�����ٌ+8x��C�)jV[������$2ۡz��A�¿+���g�� ��T�Ա5�;���h�|n+���۾ܑq��v�|�p�L=�7&4k�?1s,|��X�ԡ��(ZvP�2|CE�cq9���U�R��`b[��i�(l���GΎ�Mq&�u�h��o��=`jn਀��������k��z���?<�wM�b)+��қ�|S��� df�Q`��q�X���x$P�X�쨪�˱�x�*se;��El�ā˜i��.~�mw����
�ל�"��<�Rv���R�rQA�j�g�'Kw�eEC����\UO����5���Y���.�,���Y��v�u[6٣��vQ?�uw`6�S��?(.�|�m�l�����/��Y���=W,C(�IwJ���Y;DH�Q�1�����ۍ�;r��� +1�����������/�I|JHj��Э�z���[��Ylr������U1�,X8��$��Ϯ}L�r�4�*e�_��ܽ���y}����,"��ݤU�é�w8�?������H�5�8��i�������>Ƥ	�E�:*��)j�8|�εP��P�%�P�nA
��&2�Z���r\I���9�гȪ޵�GV��PV�ꡒ*t���t፻���L�]QU3��=���ɭ����u�#< ȁh�[����&a;OB]�
"�ԛ�Xn��V6>��O��nT}u�9��VA ���J�kM��h��p|�D�����W�����فc�}̄�	���6*�)�����
A��+�`���\��7:��ٿ6q��w�RĨ��\�l�.��)ƪ�;����k̗(ߣ�%hA���."\��cG9Kpw@��9���2ֳ��}��͖�Y���A���F0C1��]�V�y����@���[V���� Qa� �N��2 �q�'x��Pֲ� ��a�E11���R3' ��"^`��$���[��9�l��
\�5��%e�F\L/�7j�523��$��8�I� ���<���T�:�1�rY��al�2أ�g����8�Oqc�J�a[�"�����<b�Y��	�:�uՔ�͇�2��`Y��2=�k5��K;����A���&*lבȳB��lK���<a�.o��S��>�hJo���Ax/��qB�NW���5�,��H@䟩�$��~^��ָ��L�o9jT`���6U�!�zfq@j��J�a��T�sc�5W�c#6vE����?����)\�;���&����u��L��)�{t� ��(G��L#��	 U�:?��N8�>)���-VfB���}���q0���Q�i=�Z�B�,�<;�*��`5.���s^�b��'�$��mպ�u�g��wO��5u�l�ӯ�]3ά� ������g:���1#y���]#����
�c~��̟?�@b�l��#�`�fP-N�n~Y�+m�I�yp��N�!4��n��^۷j��Oʜ���[���A䷊��"F(�����HSLF����>@!����-��`a]��]E�� 