XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@W��n.6�u����)뙁g�}�]�F�ܲG�8|��Ų+�:>f}Uҁʄ�Q�	1�ǭ��U�WuSn��q�{�[�n	�ier�B�����5�PL�7�ysF}���D�|���m5K���K鰮p�SmC���N�f
f·�rkǖ�ijD�NS�BN�� )������Q�#��� ���Rk���/����%������
ā�`=��� b�����ڥ@*��g惑ȮX)�\��MѸ�J��8��}V���J.�!�;��1���K)�d�^�m�,1������ANYK�$cS�������*"u�L���cu��u~�&��"w�ʗ��ǡ̄,?V^��+��u������v��2��^8v)).'�L��.�5�R�O��H�x_� fg}����W�TQ��5�Lp"-?�"Wj�m��-��v��O�Q�Xޟ�l5�c�JkB-���^�'�^�L���vF\l@�i	6�w��$:4�}ZJ_��JA��|��sl�2���_���v�r���7�X�q]F��O&ۡ�ݭ&`���远�0����GzH9��۩�;C|lJ�=ى#Toz��C~#ma�uE�c�Ǻ�*�E�J�|kv}��j�������`���jP���H�{�(��*=z��ͮT�б2�p���A�]*:�	'�}s�7�LuЖ2%|�K1��8ʽ�ݚ*�/���ȑ�z�������v�#�q�r�ė���c��r�����K��`
i�sqI����ܿ���XlxVHYEB    fa00    2a40�3Cȵ�����;N~U�a~�b�k���
��̱��p8I)jԲ؞�d?��3�%��Et5��,�'�G�i���P�����PH���/A/�nDM��>�sA]Ԇ�����4�5t3�}�z�ټI�d쯑�_�mz?�o����>�a�{��C�t�:�M���2̪x��k�'�SEX
b�a�s�l&d�M��g�44��aH��&r��$��yɄ�r�:�\0fވ3�okQl��+C��Ѫ�blǸ��&����8�&���م�W_òM>�Y�9|���<ȓlWHbpr-��N�A�=�F�d�.3��3wWb@<�-��q��w�},�������YC!��m�;��O���m�І���DI`�r�
{ܠ_��X���]���U���:�!7� �J�Q?mb-pF.���k��ȇ5��'�Q6���"�}�M ��~儭�6�N:6�����b�l���A� $���f�^�r��;�F�-"D���,���*�Ȣ `ܩ�G���~�Ћ'n5��79Z��VKTMv�@�����_���F��؆�'���gSk�$��e�'R�8L��"5�4Wo\CS-�ailCZx��O����/�/>�'�C�����dX.�U��ݧ��+���o�m�@��o�?P؈���C-�'����^7ә���܄#'�C� N��gi����Ӛf��٠���\�,1�#֨J=��%*a���"�0}�&ډr���(�<q�����$���ua�B�f�O��`6%�,�����-��Z��S�v5[�oj
�=?!�E��XYt=�R�$�� .��"���x�U��!fgmp�Kl%�옃>�l\������/�,�M -��3�}��靟�m��	��� ��i�^[���l2�XfX�[D>l�2��#!>�G��+/�F��N[�G#e�rkr4W�ҹ��UF��~Q���.��&6�f�3X
���IWLd�d,Cҵ9�.m�����.��;?�b��|��8+�w��Tߪ��kڨ�rvٛc�N�3?�7�&�����Q��\�ǭ�G�jk�װE�P�R�ރ!D�����#����9mm���ܠ�Ͷ EOo�DC�t��g��ꥎG��lE�j��B��t�.i����)�O��P�$ˌ�v&�RP�"�/�?��i�&���\K��%���GVH<c�$LQߗ�t�㹧e��r|�.lb7��R�,����y����P�*����!Y�!�&_���hW����im��f3z/X���m� ��铩�a.�lg�]j̳���q�l̄9�|u=�ӑ�u�
��cxH��X�J�<��T��v{Q�#�t�g�_��Y�w2N9�N����D���+�
�2���'��>�쾞�|b�gt �V���|GUn'br/H��-`��GwE�D�t��� ���@�u�=�O2#Ө���{9�b~VR��@�2���j�KQ1�$�w��R��ˀ�=䑊�IC���Ϻ�"ёߊ�5-er�H� ��N `�v��e�(mR�ɬ�0�	��p���CL�vTL��ǹ��jLcb�f��-��v��e�p"�ݐ�Fa5�U�]���7���<�l�C�5�FU��Y�R�7��}-O��~_3��8���yʚIKA;���V]S�{��KFԡ��Z�����?T��-�����>�>�a�F�
�nږfv{�����Y�1y����t�a^��P�
�Ҏ`R2�<>�]����n� �C5W�H�ț���O��w�b�*@n��2s�f/��rT=)�9�։�J�Ε�&���S����� MA��Oza�|�Β�{�w�#�LD��uF�}s���Lɻ�I�}���ۏ`��3��9�����\��͊]�)��:�wVי��\ء6!{�^	ֹ8�n�E�)*7?
��ɵ�@�- %�y��}�:v�lTFB�A]�4��H�P��F�W5��I���N����N}�l�����j�b�VZclRD��NE� ��x>ǈ����% ����?Ni��Yf��w�|:n-�2d��[S�`w�k����_3���쬛iB�Fր���|ƨf�g�e��`�[�������;����Y)�ᬙӜ'*�p��!�Ip���n3j�T�I���҆>���x@��-Iޛ��k��8hG��/`��%#��{"�Z�hG>q@&��T+^�f�q:C/��$[�e <×���}j�3��k_�6��&oX��-�Fn����3϶t��gX�rxA����d�/�4���μw��d#�H1�I"%���͡�~>9�����$,�^]�;X�;��1�]�k���V���T���f�j;��z�4���"@CڞR]��D��>9ES��Z؝���+���-O|��X�?kS�!c���t�uG_i�qȼs� �S�~�{.��fs�c��0~�2��^�ؔ�_���%G_*��T�g�Y�����0�X4�eX�wV���r�r�q���?����z*�D�	��b�ƣġpc����e&���3�bq��5J������S�{��!k)�VY�p����<��t���>�xgk57!Ȏ�ҟ��5�#�5���N�)�=������@i�/���$"�W��_��;�^}~��-�7Y� �{�J��~�X7P
�SS���]��A���M�i�ƈ���j�Cw��3�Ѷ� BW@�x7����1cSG�~GNux	j��8H��`��&�Dt]G"�lG�U!�-vk���~��Bd�w1���m�="uZ�����O�-{&�3Z$ѿ�m�PaP�h��h��$ns]���'��k�00R��|���-T�+m��q�sc�֧:K�V��W�}i���T���B캰�C]�̃�D5	I��?�w6T�$��a�+�Lntvj��.i�`υ�`���z�"�vG]�Q@������vyr��&[��Î��d����'���j����F��J�h�fC�ď.�ȳ"��K��g�J���/�ه��F�0���X���`�����y����'�$��^����U�&�,��8�ְ��]$�O���c$@7��,聳�|.�B�G7�)��;�DͽۓoԵF��$U�i,��Gx�O�~�xN{[�'T�ʘ�ױR�����
�Q"�B� |��Q:��T,�����JI�zv�1���RR˂��~��L�1n	�Է3���-�p�g���>���W����k$(��!
��M�^�;���LL� bC�Y��� ��	JU���7�g�.1@��<kp^X ���}��z������6�P��[�~&a��xD�yD��n�E>�ȸ⮘,u����@��^�0��g�&�[��2�<y#� ̛�Geb�Hv��V��֐Ղ3�P�Y���͓�U
�ce4_]J}�&G?�,�W�Ͷ����3)x�i�[�[g��p������K5�����ߞ�Њg�e�����j��+��Nv3HK��}��J�ja"��k1/�!��U�*����#ר����򨃰|�k����,`Ί�v�G�6��*�:
j��1�{��'̈�H���b��L@��W� ��A�d �(35Fu%�����X.���6������!"�3��
'|��fa�5��Ny�7�7�-�K�~�����p�B��ŷ�Ӝ]�$V28���
'��s�^؎��J�w�A�7�v�$�Ps�0���+��?�؈�r�n��񮉺��.�Z�ģo��1����в�AMe�[���3�a:��빴���A�|��JTNM�R���p$���S4��Z����h5!U�+�D�2O����r(���O��1�^�F}���M�i���A�=���2Q���ۃ�R�Mp��J�R�@�d�M�
u?Dn�1��U��t��o�D�� �=�`ޚ�Ԛ>��a���γ�nϒ]Zӝ�G�dz����T�
ۗ���X�� �zߴ&���Rb�K������I p����K�������:B�Q4n
԰�$M;&��O���J��_�R+���v�<��-#��4?��u3���]^����ë���X@`�n��LjU���S_��eE�^^�1�t�J�Y�A7����wݭ$���TEz���Xm�.�(�k	R핵� ���y^
����=Ez�ܟ�8z��(�P�S@���}��z����X�n>����l�(��OLhs���
IG���C��Q��<<���	=<U����X�|� z���
MZ�+`�f�i�zl�cQ��W���{�x�Պ��&�k�8��2��i��R8���r�a��\�V��6gY����A8Հ?�b��v.}o�������Z����U�rB�]{���^-q@u��u����b��˒}�E�C�'� r<�6�ayǎ�G{v��QX��ܙv��|x���?�����bq�&l6'�pP�B9�O�},�*Ԅ�s��A�r�Xz�<�63R�U�L��m�*�:-E[�F4��?$��K5�#l�>���K[��h`%$[�ZC����
��ݠ�m���5���P��ߎP¥���C�SD;���c;	�l���Dq^�B����!/�c' R�}"�����w��#��q�Wǭ��>Y%�
��*)��'w}��*T���0��i����˂E��Qg�`��cNv^��-3������R���c���<A���X͏�;$>d��V�^���(�	DU5��8E{�mon�#��C�E�}��Ҿ����d�(�ݞ���d`��q~�Z�)��{,��Nb8�3_�bI�����D������>=���(^BVusD�ׁ��I�|�Dc���]⚍�:z�/�X�Q�DO��,�J� �X�
����r���+�J�ڢYsۨc���X����Pb�?��=M��Q���&`�a.5K| s��6�j\�����\'��q�ek���@sΏF�P�H>}����ê��ݦ�T8�!���6�|�u�h69� ~����f��2��ssV��Y�Y;MhG&�=MF��S�8��@6�N]c:��{!*~���_2o�M*!�(A6�_�>��~˩�F�}����l�!�`G>%�'*�^$ơ�Ʂ΍ 
�B�P�R����c�g�yeHF&g����s�_�ޟex^��q;P�|�r酪�L���7궒��p�]���+�����@g�ԶJ[ZI��c4.��uf3ܭ͛D���C�qqwj�]�_|��ұ�Q��Ͼ�\�^���oHS�Om�n^�U:�5ӷ�SG7e�=�� Pt��t\Qr@�9ܡ�p��>�/�3����a��~ئ-
WrJ�|�r�FfL)݁X�~ $��\�W�U�6��_O9�֎[�۹��� ��?)	V?����N�f�3=��l�VR(�n_��<U�=R�D��{b��,���l𡷁��k19"�ё���r���'���^!��f����y�\k���6&3��L�EP����թ�<���w��D�9y��.��eh��{�]q]/3�!��]� �Uo��;��&�S��	7u���c ��V���X�����{�~���K��D���4��Jڱ�	��z+����ޱ,��y��Vy<΂<k�#�3�Q�Kq�I!���
���W��ᗆ���΢�^����6�0%�KZ=��ZZr[�=[��4̥tA�ieX���N��N��E�T��a��Нm5[�4W���4J�LA+~D��WAd���)� � 9I�����d�^�g@$ώ��tGbŁش��T�(�j�	��h�~7+"���0���,©\-�Q�HG~��W�Y��-�8��륇��l~֌yC�,]dE$Bwi<D��Nŋ�T�"�88���	h�y�i�ai=8�avՓ����~���eн��}1~`k�$���P��3w.l�JI�P�r'J�J�fd�Dn&U�
Ѻ�5��s9i]G�/�����9�0�&د�+&)��Z�1L�[k�)�jF�a^�|x��1#�́�8��X�'X4e'������t8��h�w�9�"�����¬�
�Դ��d } �~��'A���v�ۛ�x�����&�RF��F�"qM$�8rV	euhM�����W��)a\��X$�o�q��Dl����m��&�%gf'a,(���wTsc]��Ԯ�2��::��Z��ɏ�%	��C;�&�n��U���"Rё�--6B��G���X���'AQ� �bv��A���)�m���un�]�'��,dy��gT�@��s�;��p�A�2�=��i��z��q��cO��.\��ve���4o8J�r�+K��[&�y��>��yc��x�L�@�m���b'w�Z��?�8�wnFT}����3;04�Q��ZT�A��y8�P�r�mb�R����o�eC6�.(�s�W���q�ΝA*��c��,[#�:(~�,�y�eWu�SJ�۝�O����W��{�O+譭��S#*��O�ᄩ�:��)L���
s�V�����	�*ʛ�n�r�2�/>��
l<��Ď�m��o����g�QJH��%�_���F�w�biI��Ә|�N/?3l�<!�o�x]�Brt��VQj2�<kf���e
�T=��WY�@_'92�5ʞEQ��X��g�mE���p>�V)�qO���g+ [��}n�������Ĵ�>�S�����I�Kq\0/f0�8B�f��7^sPtA	��V69;0��k�'�d"k�����3���N6M�k2�����M�mʔ��nD����wtW"wg�xzfzN��$w6;>���0���0lR��F�=�Y*UIh�Oz.���J4sX3L����8��;
��/*T5u)����*�mYcޭ���t��f��^:�2*��D`*eu��Y_!ٶ��e<�u��e�2�\����5Q�/���1'u
f��냵K&�d��o���D��}�8B�۠<��5|T����;?Cm}�
��G+7H�tn� �8��~$5ؾw���'ZŁ�h�̼�"}�͍8�'����>M^K����۴U� {wZ���aA.��pG���;
��B�Jm����)�B��y�"��D�e�A��y1sdD�3s��O�z�ɐ?~�x���R�{bݪl���2�����`cY�)l�ĭ.��KI��<Bb˫{w�
� �G�{�P����7r[^�y�qȯ��\��N_�J(ݟc��T�]zۇW�����kZ$�|���Y2��K��7.�{�yjP�D� g(EZb���_��clj�FG �3�
��4A�b3'�Ba!�S5��=�֙>Z��l+����hM���'OOCy\_��c�NE#��8���X��veh�o�>9h�'Pn�}�)�C�>B��N����?O�Y4�T���� =5�)�3?�kX�+�h5�$��uf9�7����H�x�K`k��L]S��?.��/2@��,WYT$2�
.(|��� $`��ꝩ����x~�Cj4ڳ;Q&;��JB-�=e���©��n��^�*-Nf}n�8�@��_�g�/ ��8 w�s��Z��4ċJ��bzx�n��D?=������!J>t�i'm�U�Bt9�!=����Tۈ�����vw��ι����5 �졙7�3	K���E�����sv�,W I���X�/��.�9�x�6S��M�ݻ[[Y;�8�$F]�(sFe��s�j�tPJ��A+�y[ Գ�gbx��$&�ߢz}�?��Q{�>u����u,~�jk ���'~�^�3tl�
���c���n���nNMv��8����'�q��?�4n���y�eP�S.�H��u�#7b�� 8Q�+}W��k^���\��q�>T��>n?��}.�y����"�$�����l�e�oB�Z�=%�2��O�,:�'�"͉V�/��RQZɾ���6��\[S�%F#c9A�w��K7�]1����xϣi .�A�̥+�M�$f\S(o���8>~��ūn_��Tn'A�wJ�].��}��NRo�����6�x���2��[�A*��-4Le��z���U5��#^�˲�-Ǟj�تI��R(�.����s㙑�$�4����4����6��HvQ��$*�P����v'�p�\4�b�9�A�*��Dtd�O��(�W�C5�ޥ}��^��φ���>'F��x2���u�oo��o��0�=�}@������tP�3E�B8�����E��E���%<&MƂU�Y�oN+376ז}d���d�軧WZi���٭�x>���X6�����h<��z1���בJX����!��E���
%���,�͵��X��U��xfYXqt�l�VZ���v�I���"�`~8�5���=>_��5������]~# 򐂝�:�) ����k���jˬ)@�\��Y�Y)N�b]K\Texj�h�����\Y, X�ڠ.��~V��@سlM2��t��� �@��٨�m3��[�J��<����!aJ�-�J)e���s���+M��%��i����ҋ��J1t�0�GN���3Y��CA1>��h����W0�|j�ߤ4�kv���LS��e4���S���g�_o�a��zNRNZ�9n��_�y���3X�N㝥rU���X��_z���B��0Y�����{�(��o���w i��[�-0�Z9-���f�O|`\E֔�!^BԶ�(��:�W�ROM.�4\���C���$-Ј��d�e��cW6O����!�9}#�Fa�h⤻��4� ���jV��>��i���}E���s��IB$�
b�*/*fFg	�����>V
W_ނ
���⥁����$�[?%z�#cH�)'F�b�x\0�J���Lh�T�;wԠ+�(��ģ����bW@n.p'�[@�_�v} ��"���S��ӹ��4]�V�ǫ�����]���}�����E�W6!�U�����bzL��.���QlFBS���&t��X�ﾏO�fa�A)��b�Lt7l�'�����h�u#�<*���W�%���q�Յl������i��~�+Yf<���M؟K?	� �mQ(�g·�� )���������x4J<y��=��W/�q"�4��<�J�S��emf����m6�ޛ��Z(��� 6v��g7*�%H���C�ߎ4W�?vr�V1>���q���6[�7�_�,�E�v���V�;7�v����[��;KV2zI�tIG"�s����-׃�����8�_������Px�6Hfr�u��De(�;�x��M�ě7���m���G>�y�	�����l(c���'�g(DD��C�ra)ؖ.�$);��>(�5�劁0������"�g��O��u��+c$ҋ�
]~�9e��|�d����D^;��fޜ�JiρX"|�{>_?l��z�8t�tt� �l���A�n^��M�x�(���W]�y�]�vBNdH�����{�������^�E�w������E��)�1����h^ĝ�Vo�Jw�S���z�5)2�H1mI�U
��÷W��z���=W�`����c���^��e8/"�*�@I�[�biؙ:�"��4LmJp��nGJ_�)��~7�ys�(X��R!jn�[=�����{�5q�f�fc!�"Օ��;Ό����up�ğ-y����gqz�ӡ1~
���*������F�x�(�_�Ӡ��]u�KW�_3�w� 5��J�7fť��{���{�O�^����"�%̋� �a�[�T�(����;�/S��(��s 6=�gLv����Nb�)�g��Ԑh��,_8����V[!����2ǩ*'�SV#����`ܚM�(��t�Ч�4��8k>�Ca�t�.�Po���wQ��{�������<�_�F'mB<*74�6#tŖ�=(RC��T\��{Č�>Q�j� �����>y#L�:�%�Ah�~�҃�`.�[����7U<�������1�I����QD�+�ͧg���'|1b�+�<;�Q���eb��H��v��w���7������0=�
�����qa�SI���_�va�26 f2�T4j�Am=g�Ӽ �F�SNj�Qs�����ϖ�$�t]�,+M�樹r}YJ��ͅ��_;���+���_.1���?8�d7R�����>����)�+��4�(�en���s����`�̺�($K�f�����]���Q����5Y�w�Μ��4	bo��j6
�^=�C[��B����|H����t�]��~;!����	S{��?��0�
�Վa��4���of�8d�o�)�7B�"b����~w�Z��$p|�>�Q#푹�SK�FS��H�Ö�Y�p��1�笴P?�}�_��j+=J�`J�b�̢�P�7߁;�\!$�=�wf��mVH��1%�$5�b��|cPgT@,ǐ��3`l#�U'8���<���7������á;}$�	Q��T�����e��
�)1�+������EDtG��&œC�Y4�0�Q�Qx+��z���F<���a����}��?�H� ������b�䐍��qnWC�Z�t�����$�o�����auU��u�)�7�hBb��V`�m��7��0���Bn���R��tt('�$gPU��(��-=XlxVHYEB    fa00     8e0��"OρG���!��q���=��duFDW��d�a���*c������_�X���5#+[ӗ� G��a� M�wY��g�_�o�n6�@h�$Rp;�b�V;�f���쬰u�=:G����]�*�!-Ã#�/�o�-��li�;x���C_Ǣ�ݦ�k_G��N;]�-� ���.��3	�F1��B���N��9{.2�t%��u�@
v-�����K<d�f�P��L- $n��0)���9����X&�M��r�u�	Žh�S��~O�;A��E#d]^{Y�'���L҂p���@����+.�Y˟���,|�uMh�C�#W)ƙma���!q��1A�z�l����{(�:t����u���+|�������M|�;�4$(8�ڼ�Dz�o�)fؘv�-�|���a�������F�ƈ۳ g�%p�[K��kt�Uk����ZHwI*T�,���X��N薥p�3�.�q�@�?�o������QhQ����`�}���8�@μ��I<��|R�����I�v(��)sԾ�ܸk�S�ca�34f��˅����9R�%�(� 2.pn���M�hԿ��ܮ�=��Ƿ�|E��#J�o��qbG@v�h����m��Q����3���wnC'C�uS�c}�I
���k�Ev�	o�ț=�Y-�E�7*>��E���X��4�t�W��[tg���� ��6�ma7'��K޴N�wM|�igcщ)U!2�%t�Z?~L `"o��9t˗2��5x�W�`���X.Bq�V��c��^�c˃!w�Zx�mm��-Y�V;P$w���r��pAd�hjeѤ�u�`��\Nz�/��P����(�b��A'���"�h����YA�Dxa{�mI|���`2R�LBM�y��	J����ŋa���6�-����,�W_|���m�O�S��D�A#7 #�j*_�<�e�ctC��p^X���Bd����O9�y�Tv�P�n�K>TW�	�k��������i1���J�H�X�j�����&�n�+�1��q��yVU��Y�[\�a{��i��S�1�Aa��V�9n����ۻ��u�����R����w��'HI؍7Fh��l0c����΀�6�!�/ةF�"&�R�U��}ȁH�H����|� �`�PW���j;�.Dn�t�(A��;u"�,�6[�7Z���ǉQ}U�H	���>H�&8�� o�ҸlzhN�9�s+����J8����+�k,�P�q�����]49!=���MFM�*0�Ź���_x7���^=IXj6�!�)�|��p�Z�@ ���:X�u1��h�����!�Q�f~��<�Mg�G����2#=��FVWah�Uf�F���\q4���(�M��8RC�(�и�o鰨�Ka0�t+L̀~/�8�b�e��o�1�˽��b|9v*�vL�d��>�67��1_����t	�t�og�6(jZ�ߎ��d� g�ōi�q^�i�z�����$�#3j�G%�%��G��s�^_��[�T���嘴Ӥf��"穑��u��ZH����˿�W+��b2��/� F-���g�������#uBC2��"�
RK�yV���2w�T���/�ʽ\s>�����Xw��0`���̷ך[d��y"� ��u0���y\.t��d(1��|~��p�@1�U%{S�[N1�`�lE:�qS�0@�@�9A�QD{x�f��- �=~|Z�l��s~-�&�ĭ��C���o�	���{��)ʠ7n�3hUSP��ӑ��م-ч�0��C���/6ҩlG������Չkz�Ke�Fىl9�Moԥ��5\�Ea�x�{]d�{�ۂ��-v�#G8�X
�j�sŷ:sd��7G��b��D����{q�$���q/��#7���E��ul;	�@�Un��#/�Ŭ����}S��ӳ�B19}ש\�8�ܰ�ה�lę�y�5�Am]�YH��ر��ǳav�t�%��cX	=YhV����d�^Y���⤕���������xZZ�Wf��֊2�tI�,Ii��������*��24� ���X��a��(����!���S��,�}��-,�a̝W�\�2�b�0�O����9���BGq�q�h���J��6�LsA�4RR~�phm�{WUl����|�s�Ʈ0Ԝ�@�&c	�m��.y(1l�¡���@K@,���N�o��q*�S9����XlxVHYEB    fa00    1110�8L�#� r<&�R@�0X��=[f���?��#�&�E�;0QOJ���w��}��FP��fiC ���v4��L%�Q�K�G��Lp�0:�ߟ�v��ܩ�t$J^#�zfwq�&�q�crs0h#����� :Ā^�tT�8��r}����Ɵ8�D�+F.�t��%��&}�	tC0��2�乷������ķ}v����>2�x*7ϊ�������L�3�W���
V�?�U��Mi��#P�q��A�u~g�7L�Q)�K�s L� 
I����@.���}�	�L.�}�"x������^S�(��l�aX?\�<�Ֆ�]�]���s�b�z��Di����r�o��VR�1�?b����.=Gȕ�A) �1�ơfQN�T:R�$Ú�G��!w�;���]῱�'��(6���\/ģ��
L�p�$Т\�����W�V���!F�!@`����d�a�h[�$�P�7��i��A�rV�2�3��M�r���5,+1�HS{��LL)�t���)�r`yj����'��&�/�k�gS.M@�Y�����Υ��
���(��%y6�4FboYD��1��P�,�;���=��)[�GKɩ��B�u�u�Ԓ;�I�	�	�ՠ��O2FK�K����OTW�R�ns�����%\��UB��	M��^�b����ĕs�O���G���g�����<�5�D2o����:��M��cy���{	���ᴸ�q'.1�*��l��m#�k;���p'B׷W��̎5�O`2Ȯ��"��3fA��JR#�zrx�w4�$Z}'
My�[�kI�E��d�*����T��WI�XVa�>^�ß�8�v��F���}#��G��#�� ����I���s�W�q֍�
����F��Ѻ�b�@Tm���ݝH�+�����=Ւ>���^X@t46v�FffCiS�:��#]����R|ap�$�, s�j%<4�`���/�	i� �bG�@�B2��=$�rt��.���^��#sW����q�_�:�/���i�ѧB�/�,��y�r*Xf$˅vgfm����0o�¢4๹�%���>>]�˵��Ϣ�a);�x	&1[j�5]x��_���u�����)���|r����M�U�A���&��"�M�i%�<�����YFnܼdyP��ݞb�b�U��)��;D}��e�O��$�c����=t���� ��!#�ڰf�����<� a���`[H�^�Z�;Vdz{tA͋��Q�;`.r��*02@��Q��`�Ж��q�/�z)B��Kj�az������!������\�������U[^�`lw^��r� �VE���c���ڄ(�OF7���]�:� ��cn��h>$XG�נ�gG���]��wz�vۅܺ��Q2���]�������;J����0���_,��ȝ(Y���E w#���&(��8�"=�W�h1��œ)�FL�N���ƪ�tk���aa����ꠞ��5��Q�[Щj!��J��$��Ƿ�J���7X��ڜ8(�ܬc�рi��#Q������y���pnpS�VMR�D��NXSN'��y1�c��^Z�;�%�B�/��:w��m�v��N]G�'��]�yF��v�`�6
J�(�R�[��O&��S�����it��5��2�۰�36�ڥ����斡��� -P�*5,�Qۼ�G�<�!e@�T2Z됴���7$X�Y֨z7TZ"�V���I�T��h@�U��1���׏�q�N���� �Q��y�d��x�)���G#�ڲ�b�C�oS����B!�il�x�Is�|\�焙��9�?Lk�c��ZR����to�{�����޲�ϝy�ʰ� ��e��vg���y=|� �f�͡Ш2�
G�(ˣ	�6@o|y�����q������Zx3�\��)GG?�zh�`�wR�Ϻ�����k����~��a���.GL���?���PS:�6��.��ult��R���運�&��U�l��rSϻy�������d���ߢ?:��,r|�!���0Rȿ;�HY�L����1�\0�&��Jv`��Y��/��1���4�&WmQ�[�RÑK3�J%u��b�G0h,�th,�i��f�)
����`Fs�	�����2�L��A�P2��W�r`��_���=�K�o��\5���+\J��~K��7�<HX����x���p�Nt��|AkY�w [�,��)���޾�*E�&4��O����n��K}\�O>&�5�>q	;�+.��s5 �I�h8J5�;� ����k�i1�VOvu��Pa-e
$��U8r��/��MJg6������,������4���RL��]�f��B� ����h::�31̗��y��o��f��Hj��ˀ���}�O1�FE9雼<<��&������a�{�ހ��)d���$V��eY]s4L�O��,��M �ֵ��?�*�us�rnQ�/�2K<� �!�R ��d2��|A{=�(��T�g�<`�u�|P-�{'mV�q1�Ŷ��*P�K^�y�1����y������E9��F���$.�����YE�7l��ļ�ɸ���治�B�P�Y�b��Ԝ��jc�^�s�Pc2�$!�Y�Xi�ko+��Qo�6���ة���M�~/�mq(�6컁�L��G��,i���WOߺ|q;����n8���* ҏZO�S�i,���nm����HU�4n�u��9g�U��&��S�ج���(���UO`�0�K�4=��s�.��S�Ӟ�p��<��
:X��x�Xf%�	ʂ����u��ďCA������T�q
ʈ��}��E�M�e�ld�<�����!��<i�Dn�(���o�*�I7,�Y��[~*zq��[��)��ɟ�6&J="�x��*��]�8B5�X��i*���.0��������\���+�kU6��&����4��}*�fxin*
��-�d�K�qn˙p�h������-n?��(���劒��Z,r[���Vo!��"~�j��-�i�
4ӷ�V�$O�o��)���5��JA3�t�t�RC��!
�����G��Y�axz�&S���0��>'���vK����Y ��0Lǆ��?���C�+#�mhI 5Фt)���A+Ұ�׀d��ܴ60=`�#�a+Z��֏�Q}��}��&�jd��s���0�1�f��W�SU,[$�9�[�/�pU���(Dbs��*��QP#�Z�C��%[��
֨)���;��yB儬^��N"����P��)"q�ve�2��A�
ԗkQ䝋J��ny�1� �p��/R �p��i��bY]@��r��E���"�4�� d���`�i��+VE���%@��,]F
�w�ΔKB,�[j����o�����0U����7D,i�F�G�km�c>w�JK̋b���4�>�߬��p��<�@��Z�ƀ/RᙱWZuiqiO�]��I�Pt7: �fζ$DEt�YQS�[����]B�qw��ҟMvV�o_�iQ�l�u!1�H���u���T1|!)Ī${��i�h����&}K�C�	˃{�%y������_|P��u�{�N11�`b�bOz��V����6���ͧ���F��wcp�,��1P�1�^�W��e�����N���e5��f��-n�Q^ۣ\�rZ$��]��G֞9甗����sb���+5v��ԄM�U�Utu^\�VW)ϴ���q��W{����P���_��/����%g$�#*;?�0|�_��^�瞧��W05_V��Ϧ_l簣�k�t�5п�;��"8~�Gx	�Q�xu��7�%I�Y�N�1q�lgT�]9�t��ڎR #���\�Hf�ȑ��]�Ӗ��/M���v�F�FQ3seN57?2"��%0S��:���8JA�h�*�A5�g��ǰDl���O�8�k�s�R'���'�.˭O�^y|��,�$��1#聙w0��1�����	5b �_/z�ߜ�]��<%���)޿�n)����=I�;�@P��'#P�c���F��ĸ1e����/���ug�w���������0[�&��r=7������!2�#������9
��\�f�:n��*�
PC��|�,N��mͯ Ҧ��LBtz�8_*���ތ&�g�pY�n�"����~U�K�C���<K�a;M��|�t�$��VU�C��RҊ��8؍��B����ŇB-vJ2�0�%z���:�y�	��T;�t娱��ϳ ;yV0b������&kWI[�8��1�����F�k@[��XlxVHYEB    fa00     ca0!�.�������#���>OϴO���H=�LV�%o�v��A�8�m��1�)+��[�eEG�/`�#����|�큜�ء����)�͋-,!޷��f��;�6 R�V��c�z�k�v���F1�~�3��Uq8ܔf'�߹;20�_�I(��$d���ھ
6k��ה��Q��>��E��5���0\��^}��?2�xk01}�;a0��o-{L����\e�)�v@��<�j�T��S�%�ڈ^on� <$:�6���Y����H�Q�oS	y��Ĝ�h ��ʕ��E7Q8�xm"ck�y��|�k�����ǝ�Z�_�-�C�#��];��\*4Sr��k��[8��-�tt�Y�2h_���N�о�(;��^E��t�/����g���	�Dŗq?�¿w��sRJ���Ѫ~"�M��à�z�#88��
����%�-	���5r�k*&/"R|u�"V&u³u�gP�+�6e!�>����˾�Q��?V�� 1���ݶ�x̪�]�w�G./{`�:]�+ߐao�Vm�ʔn�����Tz%������٧�O�Ԅw�e9[{'C�ƒ���$Ş�}��o���;��Q=bl(j<3Ik���?C�G���5o�M���� /;��X�����F~Z��~a���B.�[�T7�j�^Fܴu�{_Dhț���T�*'�ʟP:Eб��I7��y*�x|����dH��K�mA�W����&6S��j�\&%ݻ?��H�J�N�P���U��y���Q?�؃j؁�ґ#g��Ɂ��ix��-���ˢ�C�_��?��D���L�Z�ғ���:�<��P۞��H�z>~���~'����w�h���¢�7�;G�AΈ?7�8�Z�C�kܵ.�-�ua��)Q&4�.��0'n  ���.���K'��wV�(.�Ϳ�cnol���gw��髜��2�	��)��@x�� ���~x���)U	�n������J~���p�,̏��Aa�hɣG�����UW������.|�������X5-k��$���-�l� �un�s��ӴO��>3)c�L��<�U�l���u�.f��!H��=$���I�s;�A�q�WB�۸��[yr����b�^��%��(�X�'0��u�pke�ti��7d�\�u\�ƨg*5 �kP� �a�e�l�.�U���FS�� ���9W��LgK��Up�����R16 j�zf S�^�r�m�,4���+� �
�xW�a�t���/`����7��8����D�g��%�G:�� #n�F���ţí,�W���X�3��7��˯8^��6�OY���R�+��tbF�����N�Qr#���#B�0����J��`����A��M�[�H���
2gɩ�E>ٲ�g�b��z�<�V9��u� �b���C�2�DJ��c�w�#�x���5f�JͲ�c���{8}�p�^��'ʼ�Up�QS�Op_���\e_f6\H��tS��O|(N�Y�,��8DF��}�[�B��\�Y����Q�"�2���Q��U��Lq�L�W��|z�P����zkVLG����E��}�������,���1v��l4l��i=�,c�][.,uh�(��@�����@X����k��Q��ʮ��v���D�Է~��z�Ü���C3�f��9����+�A�9T^Y޴�/�y��%�x=*h�O�J���(�����ߵ���)�8�j���r%���mR/�l)�+�m(�2/�ī&�N��BdaKP?G�x�C'�=��Pl0��W�nOM'&���vW���D�����C��]��m_�'ayXc�F��� ��7TőG0���&q0�դ��"�iId��������n辀�>����r�a�{��Ԙb�-�W3o&��8�.Œ�q�F"�����W�I�,7�kJ��+F���h>>�v~���"Q���3��p�[v3�I�	ED��$���򮓡{�I?C7��!!�	�F
E��g-�^H�k�rR<�G\,�X��a}bŲ���h}ڍ�0F1��0��G�9�X�SB�AyH'l�)ev.�,� ��g�I�퐡����+K0��x�k�A��=+'�UԽHBQ
P�,�Լ�E>�'�nx�#n�/�x���4��xv��t�<a�Ez\$�نk5�I9���U=�od:���f<��T�oηe�c$�BK�CA2�{C�)^���bRh�^r"�.��H��K�#g�d����ml	�:�?m8�/��QY�2!Lq�#g"�F�[� ��f)�Z'����z-�J�� K��*s�(�FH��z.nޮz��)U�r�}%u�*��#�3�o�MU4RR#���I�>�UF�Ō�>���\�� ƠemF����ɒr�Zj ���|[$��U&E���P�� ���v��A0�'�n�=�����
�g-�	���qB_~��S�|{�Ww�i7s7�5w�^�N�c�W
��u
���(%ɵe0�3-�KԡŠJ�۳����@A#Js��2�={Xx�)�^SQ�����!X�}��rk�'�vW_ԮS./5�R�d�����J�M��H��"�9�0^��m!���H�~�B.�w��֓�@�k��/>_O�d+��Pt�.K���4Oz.�:
H*�&笧q�A���i�5�d��͖8��5s~�>⏌!D	=���s���q���P��Y�.")"^F�2\R�C�������D�čу��V	�����|���Q'� S����$}�<�� �=�c�une�4yal
i�<�l��
+���"�}���fJ ��c��A�8�L&�_���曕!�����R���*L�U���pS_�3{�+X谇?H	���h�h�Ҝ�)��֬�c�0�0&kZ�8WV�u=�%w
��{	?U5�Hl�i�w�L��z��oI������2)���K����k�v|T�հѳ&�[�^C���.ږ��2;`������c���/1S:e��q�М�� �b�-�����o@4�>�R!�ȧ���U�� ׺�x�X��{�ʤ��V,?�q��]j�����j9���׬d/-�^
��)�H�f�d]/.j��UG�kG��Ut�B����Ɔ]^��+<���c��O��]�=�� �`��`�ry�\eT8Lo+lo�4�g2�Kz�"4�GGN�����*G�_��9��j�c([��a�9�'�XlxVHYEB    fa00     3f0?���BK���>��}n<�&`���[h����莇����0tÝ��f)2ӏ\��.�Waq�p��U�k���D�;x���s�0�C��#����־Xo���V��96��[O6��
�ȌJ�{cq�>������m8��^g��X\�dr:�4/��f]r�Mfs�J�/�xu���;�3�O��>�çK�3b�~�|�Fm-�J/G����xI�}�h�������$H���4jP�qY]wc��9h�}��}��f|<�A�ʮ��5a��:C^�!7��3x5���Bt���g�v�ȫT��o�*(��+ۖ�y���c�e�Z����- vB�/�A���{�^�� !L^�(�5zvs$"��գ\�wa���/�NzU���e��p�������D�C�s��j��eiaү��{��U֬�竻e7V���]{�W��FѰ�;Bs��[K�F��G�;����b�Ⱥ�cM$� �6�r.��P��K�%ƐUu��2��%Y�g�@��k9?��9!!��!�Vw{Խ]�7POW���8�K\��1��o#�62�l�yLl����}�S1�����q��V|���)1�ωvj�["���P���x���K�uN+'u�w��1P&��Į.�P�o�ဦ_*3��Cֱ�Twԇ+n��L�PeЊ�w��х�q�qB��N��RC�`�q�G���Կ\��HC�4��b���R�N���F�BY�~�m�&���/~#�6|�т��̴an�-ro2O�mQ;�h��?��r���J�#g^j
jq���;�cd�H���&�k'��x(}8��M$�o�3?�餩0f%�2��J/��>��$�����G��ʻv�<!y�W�FK��[�/R������ԝ��^C�D�Oyu��&钼���61R����-x��d�Br����lG��W4ϙ���������Q=~FzՓ�� (�;�"�\��u�E��K������0l��$掦����4
XlxVHYEB    8096     b20>�ԇ#�2`�?��!I����ݮ�A.<P�\�������ݐ�S����)���?R���@�ș�0�y`���M�ۼ�3M.=V1���Fx��v �`��i�}|��z���x3�<��с�ѧ�S��I0D��	�s��"���a�`��k�pZc%|RQf>�-�n�������流��C�d_��15&��d�S<�(�lϜ��PǴFzznB6Wc�h�ճ}~��-"U�#���-�Җ�A=aP�Ձ�-�U�Zݳ�X��P�U�l�y�[��߬�H%�Ѳ���
v#�-����I=�k��_����h��_*O�����wHM����;�a�����FR�[��Z-.0&9wH`����DJJ�W�3��J��HrLW�@c?FxT՚]7K6FK���g�s5f	��tn�`����A���3���v{^@���YυB�)�B�*�=��4Xm�c+�g.�<۱5�H?���S���,B�nE��*H#�����A����9�㞄���
w.uGl4��X�.X�Ƃ�����)�B���ZVLb�%z*��ţ��7�k�Đ}8�O�����V{A�c|�uhgA�3s7}���u��T�\m5�gH���!��d��L� �F�!�G�4��ȕ�E���8�0�*	��<-q1��������V��kV���"���8��|�/��J�-H���4�@_L��(eؠ%9�}�o�Ǚ�ԥ�R_}���e� �F��L�H���b��խe�:�ՠ	jt�b��3!��0o�(�>@���q�(�/���Uk���nN�AN��{N��]���Z~�}�p��x�e)�d8�09����ޛc2�UC�}4��#���et_	�YvhTzn�AF�����	`'HL�O'ᮥ��_��,��_~b��f�g����{�1l�ۏ�ZϞ;��vQ¯֍H�č��ڀ�f����h�݅����M���,��T�0�Zy�(f��[~�A�s��yꢞ��xSrZ���@ rI@y�j9Mv���m��XU�����Ԏ���w %���<{��@�v��ml�|��6�ka�B�
��4tZNN.���[R��(s)�`��A蚿��ؠ��_T�j������b��e��s���a4i��I�u�$S���9�;���07�CL�<�fJ��)$C��g4���}��L��2u��`wlz�x�7O� Nj:�ӥ���u2
mqj������Q_�ȱ�Q�l���q�U`�`,.dfN�� ��G�pE�/�G-���#���b����<������G��P�YR�jї�}� W���tj�K30�Y�}oN�K��Q����7��lw��3�w�/��L* }�a� F��Ε��
�~�P���Z�@��_w7�/�WA�J�M	0R]�W1����0�۶�Iw0gx��Q�	b1�a:���\�����c��cN�v�`�Bv|PAI;?�S|��aC�xdf�� �'�׬;�Tu[?|���qL�[��zR��F�t�=�DIr���,ڽ`ǈ���\)"��N/TkC7���������5fF��$�?� �qbq��rH]4D�PDǓ����T�2��|��]y�썽�k�dv'�D� �h�a\����X��0�I��N�5��c�U�WkJ��v�7�2�}����@��p�����Q�5���OLJ�{�L*�(�-4H�l�E$�����*9���HW�0�pp�*&����3~��O@7���Ժj9��P���	&������iF[�!Y q.���dP�zE��9�)����H���幔�cCZ�c;<i/is�s���}Y�Y��6)��4�As��ɰ-3�g�؃�0�� �jJ��F�4@^i�_:Cuv	t� ��j����v�l�%����.͢o\,���#��e�C�DPcEl&UUWB�\�/�\��B .�"�y&1d螢A'�@I��{�>:k�����N���7z�6�M�����*��b.���D�wDٸ�x���u��� y������r�A�-�p������d��I٤ݯ����\g��نizJO�3А��=)�<){|.���2[���*n&�<�
H������o�F�",>Т��@���,��u�푦q�e�'U��Q�#�޴�Z2{���SV�\�Af��-����Ο ^�vJ�]��ow$$�8H�'g��;��q��*g?0�ωSh)��q_�h"�)�{9�2G��₋w�pg��*ɘ㋢�!.K��H�<-�\�6�3�mq��ib&�<abC�Q� ��D�E�tQ���?-��ao�d�8�Ct��p<����x�'�����:8�����F�K��?b�Ɲ8�^7&x�	��s���e�k�3:����^�B�5U� ]Xu��9�E"�$.�n	�e9�_�#m��_>|L��L�
�YP�9|[�x�������P��!P ���xL��I��X�Ę�<�^l�Yng�wZsb����h*XV0�h c�Z�_J�lw�F�Rq,Uݮ���IT��I��&O�1r���^J�Z�/�)GCƪ�d"����^Qc��7ZȞ�cD<�T��<+�/�NT ���dF}�����h'M
��.TO��h~gh�zeu:�����z�T|�ӹ�1�7e�^V����5�:�z���lz��Έ(TD
�)~�y5�`�,��+�XK�z�Կ�Sw�G��;�]f�k�C�V���=��#�v-x$�(���|��Xj��,O_m�b'�A��xǺ���r�x�6�-��pI`r�x�X���螹���h���