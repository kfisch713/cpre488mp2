XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{k<��ƞ��^�+xw����UIbUq��~�F��}-��� ED�U'
���#P=����k9ģ X�o.�������?D�ZH�|�!Q`-u���z�}QEh����K�D��Y�&.Xp��תvbmi�SS�Tl�C��<�ca��Us��7`0�\�����w|�봡@�Wh����Z����	K�ɮ
Fv��*��N��:��|P��q��ϕ�6�ܸH�4��3��q  �9�$"2��9k�Hfm��}~�յ�c��h�|Q��b�ݦ�Z��cH 3�E��U�l�����)%9?���#2����ʫ@*����]�f -2�>�Òp}K}���I����M�4�S��+�W#6�fl����$��E+��ˬ��@>��L�~哐];�@4lf����S���a��' ��U���2�H=7-�>B���8Y�:J�~��W|&�S��[q�l�i+�$9�ts�.��࿣1	�_c��6����uP^�qB؞+�/*@e=p6�^0�TDB��*^B�q,N	]I1d)���"b֖iZ�:4f�<��L�����$�}��f��>�*�7��lXϞK�ej�j(K`�8�Q�� gQ
#Yp)�k>��8��*&�a%�٢&.��n��P�W�O
���Q.�ln���.�����U����$ ���3	ڣ��:|�!�RLs��CN��%X�x4K+�{�z{ܱ�Ќt��.�?�&FfX�7��䎕�ڕi�;��N�����WC����"���iq3u����XlxVHYEB    3d1e     fa0\Ɇ�8C��>�?NK����.5���ર�dϾ.o4o��W�N/�T�|��6��^��������=sS���6J��Q�=r�c��c&�ƨ����]�ˌP�"�����OL`�� T����z����J<dPc�7�p�Vr�54#��Y���\�ܾ��pt�jR
c[S:3L�\��U����_jNms2~��!Q��*����R�	G��w�K�0��_Ts(�'�_�{x�O�%�D��Z�����5����J�MS�9�wS<�>A�8���f)��J��|ғ���i`17���1"�?v1�)$wL����x�(�`�Y��	,:S1]��ݹˆ��,�%�[D�r.&��r�t��}➎�M55��x4eE��9����ƻF���a�N�����5A���W��pgN;J]��<�3܇̛y��EfŜb��c��|��m���kqs���QlC�ɚ��[�hǲ��#�v�ڹ��u��6�p+K���p�Y)#����@�K��WLK� z.>�����0�m�|
��C+2��ck�4޶ ؃��p2b�@��3��;�e��C"�=�,�9S�Gh�8\�5�\0�z�OobؽF����5�V� ϩ�,fD�ƺ�f:u=�O�)���	q���l�`�s�ŵ>`p���,�p�  .�}hT��8SiA@�>�gy�>�?Ϝٱ�����ߺ�s���)�M�s�!ػ4��S���jt��J��[ �\��r�*.��	�k_\�ib�ܻlm�]�ϫ�˶e�>�e�_$M;�;n����۔1�]}ǲ��7��i�/t�]�(��4�$��������s�G.�Х��1���Z6�s����B;�٪�D����(���9���t
���+���������2�W�������0Q���T��j��} 6��$]�G0e��ϼ�~�b�WfMI�p�H{��8BEl/t�q��&����͍/M��<E�+��z��+�7�����)"�T�I����&��(_
��|/h��k�A�(I���M��`4����G=���\���-��5���YMi�K������-Q��ٺ�,șvd��~m�����2u���r$������f�����e!����-��J�;t�q�'D!`	�#T������c���l�ZC��az~�w�H�8�L�*�~[N���z�-�T���_'��pp3rC\F��~�N	�Zs�'S,:^�+:��/�gL<[X� �4�>(�����6������W��$A�c�H�d(��m·;�5�a�F�}�oG�a[�H�}K��_�'�tn���4��8��������5���wg���)e���R:e��Cu�E��+33��d@deW�7�Z-1���ɜ��G��>>�B��B2os;�{���I��Ǝ�]�o�!��G�NIkM(m�A�`�3�޾ɒh�#�U	P��Y7v<N Ū��"�H����w����.����<��S	���ǧ�1���ע���:4j�ĳ�)\\JVjxR�\C���9q-,�z~S$��z���o�9�(<�\�X~IR*��,���ށi?/X��tp&/B̛�|4��&����A00�X�`J_1��2�)i� ���;W�ǝ�U���(�i>Q�V���M��;��z�t�R���A����Ҵ�yrܢ^T�G�$���0� ���eEg�}夣D�5zu�K�G����E|��*f-ð��w\z�ci8�����*��QIe��Z��,���ؕ��3ȟ��<G]a��4w�
մJ���e«�<��'0���U��|s.C*�,��u�������SPa���X����&�.WD�Ϋ�;7=��jFr�k�U��B�����:,X�F�ٖ*�d[��i"=?�m��`��k�K�ߓ�2�Ik�b�ʕ�}��wd���'6����X��n*~g�����|#�^\x�7R/�ĥnP�!!��9�4)%�Y�Ӹ����!��?��ʍVE3���b1y����=���cQ>����[�;h��E@��˧n��h9�-����9c��`	<<�$� �I/h��N�K��o���\�S�l����P��`�C��h���	��9�)�q�e!��a�ꎗs:qU`�(�tf��k�J�V^{N:�BO�o fXqҿ����XS�Y_�Y�9L�(����C��ě��#sA��
��6zZ�c��4-��}:�5��M��Z�#z�Խ�=,`�a��u�׬�T�/�N�O���d�5�v,b����^����D\rd��ױ�ʢ�G���̀��p�E:H	H���j�Y]e&���*�GT��&�,/S�2���i�Sr$�״��3�z0���'��F����4��l����;�wb�}�������{���c����f�$]̧m�|�rE0�>e�2�=������i��nd�Z��2���D�ŵ�e����U�H{>23��R�/�g�6~!*u"��ڷ������!wa�X�M�Z}|������k�-��:�ql{�>7Ɉ�$-�P:��Jo���x{8f����%���h��ٚ��Yt"+g��'̪��������_�M�a���@ȍL���!
����g� �|��.!8XE�D��v��s4��D!�r40��=Q�*���a盧�[.6, &��}݆!ݐp�<)ʩ�\������W��\���x@5�f�	��!���� �Y&����	��0�ˍ��A�]դ���D���o���"�g ?�M��*w�C�m�DR��`v���(�^şEuI=Lsm��Ǿr8A&h2�D�`�Q���167���UDt������~���uI��R��ˎ����~�T�ܶܶ��TU�ɒ(0�x�4��`�V�e��EX*�љ�Z�澠(��A.��Ro�r�1Ql�O����Ձ2���.�~_�x"qP	k��6��k����Kk��?��TB԰0���)nd^��u�D��m�6����-��14���F�N�Ǆ��!��{�
���x�7�z&��Q�J8$���.O��8Α���ı-Hܴ��tE��2s��~M�G!|mN�/i[�':e�k�ޮ��U��$D���/---����z]a����w��#1�R�D<�J1�m8	��X��l~�&#�[�J�I��Z�0�����<��2ί#M��s|�g?��v����)͇��@?!��V/ ���L:�S�'�֢e��y�Erмu�I9��5x��,q27�Z&�E �o*��:��R4?꛷\�n��[WU���(v��4�Cm��.���c)&���P�I��F�g���P�]En=!����ʠ�<P�lb�=��G0�d�\;�4��P�`���'�L�/ ��K���c��Pq�+���Kt	~�3݃^u�����l.�N.j�R�k�mK+�3�X����ќ�Am�+fk����	EFP)+��g]5 �5d��CMI�� �iD���tX.����!���]���%���E���ΊO#��o��4�#l~�W�/s��������Tm�xR2�h�Q]���]��>U����tK�Y)ӥʊ^l[]���K5z7��a��jV=e�ڌt6��))����	㵌s F���><���Y��
��}.p�?a*��3M^�}��G�~��v��|h�����k�=������;�~��C7
����Ք�o����?]S�V�I�k��q&��|�s��Yy�9}���>A�BG� ;��,�`X̯ak/�q��]#<u��;�Y��5ዌg�}�Ŭ�V�����sL+w��Ջ���y�#�g_$l�
���?�n���B�8��L���`i��Ψ����J��A��i����y��$���