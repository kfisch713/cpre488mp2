XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��jeU�Ps�W��}�����F?'�B�Qt5UI���bY��Hˢ@aZ�1b�$7ξ���f�뤺��\g�͵هt�L�E�-eǶ1%�����h-���0	�X)rxc]K�c���k�B��)��L���4ψ�}R�(?!�&�T��?9u�i�K����w񜶦v��+��xcɍ�t�$�됝��zS�c|~���}"4���]�����a�vY��� ���{�Ǔ�ޙY�לI��@B��^���A�&� ��;4Χ'��8��\�C9���\p����bZ��_��{���B���	D�`�5����y6íܒ�Ӓ��U_�ġ�$������
2<E�g��K0O���'����":vfӪ��C7;S~�T�t3�>[� $E~���tUy����`M�D�e��^�U�?�sK�O'D�g\馟�c���R|�������Y��	��@�Cu��_0�
��L�͘�YJ^�aqF�Z��{��D��V+����P�	^��C���}��>ƾ�]�=� �ȉy�5�=�'t�⶗���gM�K���r�_��<���4�z���u<��ѡ%��z
O=�xh�NYc��6�ٿ��&H�B�b	�j���J7o˒V��+���E�cj�J�l��ρ
Q��`���>��u��_��v��g�Z��Ό"$��;�t֠���zȟ�L�1��0z=R�'.�|T05��!*��������^;9��������]<�_���|^`x¨AuXlxVHYEB    dd8f    2160�]�k|JX�=��1�?c�`�������#��l)�����y��;��I<����e
3����E�AtpO�|�]7γ5�Z�1z�&�f�w�(ycz�8Z�
����f�G�0����9��0*�L�b��σ�I$oƧu�����|݉-#[U:JD���ŏ2w�x�[�C��4��V�k��C�GO{	W���Z����F�>���d�NeYYOh*�\�j<�[��S�\$�+�9���J�D�y�Ћ���s�̻:ֶ�*���]���+��(,�B�0OA:ط
D͈�YkO��lɸU���V�1�B���в\��P������r�m���L�A��;ʫ�,d@i)6c�ZR�[��������M��?f&t��&I*�S��ƌ7�ןY��1!8i�ŬCF��D4(���2��La�������H*j0P#?x9�v�%u�F�+�;��.�4���<�%�a4����:!Aqk�>ųD��SZc�A���-G}6aU=
é�����5b"��4,�r�~��%B�s =k<�JW�'�~ h��T�s#����{D���A���&�:]��i��uZe�B]Q)oGl i�!`�`*�/�b	��+�/�����p�5�D|:���RX���iZ����^| 6��$�U�������u����ʸ�'a|�+;�"!�T��7��:�M�U����O0չOv��p��(V�	�(�=$H�1�G�`��
�F"
^w�{M�4�@�7aї�G�|L��	�S�a��CYZ�%�a���/��&�Y�]���P��j~�Ɍ���A��!*�ИMN� �p�P�@��'��eAf�P���+1w��F�gY���4xKqju1^��s�!�>A؅qZz��m�M�k��޹X�Fi(�3TR�S��Li����2��p3փO�u�恜�+���F���M�����u̴������ގG���>��hr���aV_$�����{Pj�ҠY���9�S�����ƲLX��9\9-�(�1��H#�.��t!/,�l�@���re�AR�t�ŷi�e����Ţ�ae��3�4s��KDsL�C�J��D^����{����8��o��vJ���Oy-HpS��e���
�����o�,L�՞���Ix���JJ��
���H企�m6��B#�kV���p�?*�"��Dx��E6�q���b��I+B0^�	�,'��y֖;�ة�e"������/<)�4z��x����@-f���!�9��E*J4�L�im�����Du���,���wk�ܜB��yT-��G��G�	ªMv6������uk�p1c�g�(�Q+*A-�_ B+R?񈯲�+29Q� ͍;��AS�#��=�E���$R-_��ѭ�{g�X���%�����Fn��6E�������u=�4��ugS3������}�r�.���'�ʽnDD#�b�w��;B��b�~wZ0(_�a~!���V�*���|ݲ~q��t��1rI�z(��S����.2�N�'�g03�؅�^M%����]|lR��Ղ��t���l��.+���|cj�G?�1��R�	X��C��t��O
�N$pPg�3b�X���Rf]��Ƨ��|�r�0�\�R�(/�?Y�d��ml�@w�1����/1-T!O����g���m��sQ���Ť��Y��s�{c$���K*�t �G�fp)���.���07Lb���B����i����0n��	4��p���D����Ne�=�%aLr���v�dnS*W�Zɞy\dH�F1�h�p�E�N�IM
��?�=k��Tr.nk�A�iR	�2��?�Sgs�(�J����B����B�K��vn��9�Sr5W�7����o�T��!&�K�E�v|(����o������JY$,�fp�L��@R�����S7��x=�6q1�=3l�I3�J�Rpxv8����4���%w�ށlW�1�7�����o.^�ݕ�˜���.Y�E �JS��4����?&[ך��>��"b���ͭz�z��wع�Î¿/��IB�UX����m�HWA���U�Ƣk�ƥ�O�stW6�/��߅-���-rn�J�W�i>��bp�X��m�k�1��	&r<i;�;,���:7=A{`I��Z��f�%Rɣ�����5�C<�gEB~Z���P.K�xfrT�䯒pF���̰�t���C#BIPK[ɣt1G�-�������z�]�]��z�8��q6��[��j�>Uɘ*B������s�.�|��B��?��N�������\IS�����ir�EX��y�'}Jt��mY�溌�fw�bz��^�� ��W]
��q��h/��6�i"��"�_ͽ"����t%~�ONf����KpV��1ٝH����,�R!A0��H<��������t4�'Jz;�2Q����	�e�r�SBK���2n32w�� ��A��C֭�RO޲Zf�x�%u}���v�ѿ�(�B�����*h^x��6_Y	 �VU���E�5��3+;i
��n�*�?aIBW�[��x]|%��9�"�\PU�{��B���V���T<� �έ;�1P?'�?��H�:*m�`g�2c�ɎT��Z�qA_���F+d�o�R87i��b����a��3�V�~�鄹�[�C�'���Wl��&@���n*��J���+ā`Ђ�N��5fԓ0!Z��G��Z\���_ѡ݊�=�U��a����zf����c���D �^�@�RzZ��g<�e���D�b��X6��ot�z��ٙ�4��ʐ5�&( s���f>�"��R��Z=��U_`���������"�[���؇�vF�ph�Á��u�RH�K-bч�i0��zْ~�iW�v��m���X� �$�G�KM������#�f����y�z�[���0���p�K0����X�;(�Z<LO5k����������o6@<�I��k���9M�F	J��>�J
 Tm��%ol���*��zGY7����
��Uq\�}�6��+¯Ē&N�4�w�f'��h��Z^lq�x�
E����n�=�tz͸3f�)B:S��[.ϳ>�{��9�OY�l�6m3�+IN)�D[�p1����M�n �r�?�5@��r��:et��>��w��٘S�W��X��f���Ƭ*�*��cg@#1$6_����r
��x���x)ZՌf��b���N�z�t1�E;�{�����RB`X6�)�[jB �3_`b�r+��?���l�A��f)�뢕)������ ����y�!��D#�e)������R�h��I�,V�n+|$��rIJIH�Y��W������qϿ� c]�	_K��Ǳ�ڳ���f,���<�>ש̄�͛��� ��M1���^�}+��;�Wޖ�vt6Ƞ�#bV�ٚ.a���mk��B��g$��{lXF-iFƍu�N,#c�>%�EU"β�N8�e=�fkV�������|n-.6[�N_o�'|EM(�DsCU�E+&�]�9r����MhQ͉�����/�@�Ry��<��1��|�4Z���4!���^7��z�.2V�x{�?�z%^<.�Ms�t���o�'��H���)hxHJ%nOڎs3"uꁶ�0��	���	��lZ������A���v��V���J�M��{MZ�0��<;�bzQ|���<˵\��3X~��ag�t�5��*;��O�8��8�'�N�����o|4#Y�ƭ�mV�y'��ťV.���Eh�/x�i�w�D9�o)��#~z	 c;�=�7�^���ͬKz�%�m��j�b�D�����y�F��bo�����|$���f^Dk�L_	�A����'
Ce�]1dc�k��P��N�ܳc�k�]zl��NV[Yb�?7�?��Yy"p-8J"��7m�������r��&�GU��Z"�W�8zZ�I0�L�@�Cԙ\�A�8X��VҪG�P��x�7��ú����	�<,��t�⵱9�_�=X��{�G���T��u��������f�� ��b���=����5��z����G~Z�(St�G��gʲ���q�;���H��Dq��;�gd�Q����;_�`&����M5�]L���X2"f��[�V�
��c�	��"�@�Ϋ��I���}"͵�~�j>BW�3��D:��n�0C�)Al1�A)����EEH�[�W�L,�������7ƙ��e���,�D��F���f�Ϭ�K�rX�{�{���H��0B����RZ��)�j��'.�{; X�(��K�@¼5�VV�r�����l��~O*-´�؀g�֟T�$�X�چ?P:X�'�����3�z�4	�F������W�Ȓ�3k�|0�ʤ���@�ߒ�ߨN�/�h�5hrX�*�R��n�Wx�W�R>a�J��|A���\L�i�����~$ϋ��h.���S�w��$2��AJe)%V����Xl������p'I�}K3O�7��"U���}<Џ����'���3ع �'(���$�iAy�S��f<* Us�=�������1L��)����3T9c���=eRAu�E|��F7��f�a���hm%SB?^�_��x� �JP��(l'+�^k�f�� )d$s��f���g��'��Ќ*��Ns�sBY��[H��E�zK�����e啪xQkuV�ם^��ⷣeٙ�m~�Ε/�ɒ���6rszPZ�1x*����s-�����X��2�>�\<y�j�C����H�������ߘ�8"���.�+�硒����Wz$}��?������X2��Ŷ�/=��?m"g���~T���Z�������5ċM�4p�|uKD�©�Ab:S4�7+�+P\��%������j1��`Msm�)Lu1@\�����vF��/�Q#S�o4�VǝNs���Z5le���o)�dZ�NdftA�+����Ԑeav�@ʨ��[�ؠ��S,�fw�p������LD�����]��tYB�(t(s\h�l�s�#�j7.��&c>=��K��Wl���FLq���֠�h���:I�L|q*	*
�=|iZխ��K�k>Zg����;"��\��'
1э��뛛�z��͉/�f�cCN7�_��r�v��3ZXǢ�!��tFJ#���A2�^��Ypy)/���6�\��]q)�����.����}X�Qe��L2�I�E��scns՜o����xnz5иlO��%�ӓ^�ګ@]:�&߿d:�>��PZ��ͻk�m�<�p够��Ȭ��0uEd��n�=�Y�P���|�n��_6�n`2��	���tt��*��&cc>Z�� �Xp���Q�K���,<<�M{��I���n] >���-ƛ4�x�n$A̲6XmTh���w�[/x��a��@���� ��H+��W�q��b���1�:rQS����Y��H�Z�Hr�b1	�j�:	���*��X��X��Zƶ�IO}=8+O�_��q��G�A�w�=Ձ(]{Џ�;|����?��q<�l�v�u��蛶3����^�U�߬������.���x�K]ɜ<*JM^rH�:-_ڣ�5��Ĺ�ͦ��-���џH�&���[��t7�1N+��8��q?��b�M�OK!���N�EՏ<��nf��a��n��YE�q-~9�*x��I�)�>S���� 5 �s%�.�#����
9�'��)e'�����^+���ço�<����S�=���V��S��&J"a<�~wv  ��ݓ�z|�U�0��C���Eܕ��n�9�
-�ba%�[��7�7x`d1�U3�	rlܸ�5k�'�V}��:�?���&��H������D�u�����_He۳��q�w��څv�x�Z�Y��~�2`�����V�'q��,쥟DԳ3dW��$I9C#F����]V�A�����bU����y�Ĥ�	h�h�{��^���w�_�(���*��fiŊ$.���z@��:�>�h��U�.���Z���A�@k!йj���Ԗ1#�%���$ƿi|xU1�<ɾRc�k����(�V��:��߯�aͭ!��K��.��fLj�o'}����ɮ��]#G�>5�ag?�⹛EDC#��eo�����{Y���I%?~xf��7�K4nY��
��O����n0�>��k��L������p�)3�'�A�<��󃄣`g����_�DhW
Y0?�Ds���BI!aE�G��4������dq��J�fh�2`�ctxz��|H1>J�f��d�����=�/�u�0�䥪��%U�
��1_X�톺�c�G����!��/bW��npRf�i��t؏�48�R��s�V�m��hԀb�'
G��Zy9ʼ�y"�\UFb�)�M+��]ۑ���j�1�}�(��+U�Wq��
�WR��@�5Oa(d�4$P쑑�
�f���l���\j�	k�����F�ƔNh6��v�w-Y�Tf�%�~���<�W�=�EӆS��Yy�.�k���C�ߏ�[ЗQ�tRU?jn�͒Bz���t������o^�9���9��H����i)�}��L)'�R_SIQ�#�g�"0/�MHPЯ�U�0J ^��r��M�|3TZ��b�>�8R>v��'q�]�-��M�FL�7ԝ3����?��c�E�@��`�m�0m����F��6W9Xx�r�r�yA[0.�ͼ�b����#��ن3h�����͐��6���X_�CͰ��,dw�	�2�p�sMj�|'%�|k�[s�_�Za�;�����*�ϻ���c�˷�c��xG_&Q���ۺWt�z�%>���P��m�0���9]I�ݺd�2;S�U���'��fmcp���n�e��ҍ��z��'*�2�W�U{y*U.�q�k���<lS�Ʌ�UγC�\�J�3l�P�E5L�����ß�!`ѝ������G&��fM���
��1�
L��TԎ���]U�� �B��Bc�-ӭ�Zl�*���%�;�Uj�ʒ��w���V�S��zWJ��#�n�{ސ�q2.����:��+h�,�f�h��uhm�S_>T�֗�8e0U�7���G��4q��o���:N[E�NS��Ś��鴹248�Ωg�N(/-?OZ��˖���J`G�c�\%`��)_>(_q�/\E}�Oŵ�j\��9D�!?�{��#�
g �υ[ջ��M[�� Kx�K{���Sj{$�����SG����9�˖���q7�^ܤ��10��\�Fք+�c��Z�O=���2���R�H�̄i��ME�T�:���hW.��H�)x �ً�7k�a�����Q����HA�Q	����ě
�82Q3�1�8S����aӉk[���4���U�9�p��w`��\��4�L�|��aA�d^��`��C�6̒L��Ý|=�kI��O%�'`��O�=�O.,O��v� Rz�����L?��k��{w(`%�ݨ����J����x�ȑ6F)M��mv�N�$��F5:(J���<ٞ�Wl���c��i�����4E������k(�V��b��9�
q��~��	�3��=|6�Xw{>�\*e4�#J�SI�,��5d�4�r(��C6mR;YN��a\�QŤ#�R�顩��,�R	sZ
_�W�`�o�a������p[y���٠N��.KuR�����U����V��H�:=5����"��p����E��S_;W0��"�����ƚEȢ�7g�[�sR�
�����9#���1��-�wA|D�hɥ�(�-6��<l��t_,r����8m���:����V�Ю�Ĕ�C��er|����Jhû��ۉ�4��ȶ"�8�+����l��k/�vQ{{��-�ãۈ��"}Py���`o���/��������ٌo2܄#��!�h���y�G��x�wo�G�S��%�FPca�t�U�1���W/��*��3�z%���M�:���1��DN�!,�zt�`��� ?����N���e�qoIW�H�,��_h~5rgi�O�ש��2}�Ӽ|F��w�P���¡�|�&H�bG��B��pLc����T܋_�� � �"��!u��Y�Q����X۫fH{yv<�	ģb\���~&Ζ��{��|U�����=�y�V#S���BV 1��o�7E]t�����(�Ԋ�tY/|-��=�c}B�n8K��Va\��� �#�'�,Ԭ���!ħ�^Ѽ�%�oa�f�"��h��I�@�I:<wg`�ݑ��.	����D��g0+S��R�u>o���z�U8��:�V��4�@P�0M�|�� <� ����a�M�ܦ����8�ս�ϼ�̕$��h��~4�9V/E���2L��P�d(�57�$o.��3[�~10�[og�B<>8�
}�d&���C��v�?9g�������^��8�mE�Ʌ�!��6u��8�tI~cWTCZl��Ӓ��]W��2,;�F��(+�