XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���2��b�����+�A����nq�+�� 1��ſ����B�z��m�w@;�z_�b.T���]�4S��?q)���Q;�~fG���+���[֪��^��� �>U�puz�ĽJ��&�����f	���ǘ�`��UZR�M%��� \���W�¢����gvNg �z��?�?*�/}�s�K���1y�ဴ��503k�6 ���'?�K���t[IX�U;=u	��r�E��n�ۿ���Rv\��Or��c��|� ���{�eo1X�S��d�F\J�{X�U�Nu���/�/*�"��	v�����4W�Ĥ�)�d���(��x�C+@m��1���o��Z�YEg"�`ׇW���g�T;����TC�+�UH���� ��^'���]Gc��ߦb̕c1))u�!F,���"˫*�f�%���tOiH��p��w+��_:o���N04����~�ն���j2m�g#q� �WK��b3���(|��H�U�0��	�c��Qȫn������۟�f�/F�j>�*Q�M��V��
N޳2�� C��T[�iCͬrn���]�]d��B�x�F���2��6#�[T8���!�@�S8_��
w��4tOJ�/�����!3��j�[�܌s�M�֮n:�&��"�!� �i���M�3�n���'�`zx+]}����[��w��v�>�i򙂤��:l�����=t�Z�/�"�)93����"��?�(�) �9�в.�=���n�Q iN�V���u��WH�XlxVHYEB    3d1e     fa0�Da��e_џ8����o���3�l�nCj˞1�7��r2*8�s�G�R��s���߇�����D�=�3��`��7���⻕�;zj��Ќ��0��I���q.o���"_�Y]â2�T�O&Uz'�uaC=��5PE��p�>�55R*�W��Ń�CAgěib!����C�OPk�͕�#�f���>�B��U�L�nǂ`dxT�~}XG�r��f� �����͎��~\⮨�ɀ�ܜ2%���"�)L|�����1�@�1d��u��y�ܓ>��w��'p��`;��k���o���HqP�{�$�n�V쿧���c/�n�ц��΅@ɔ��@�N��4Qc��lBQ3��;���n���J�v�vJ�#.�\'J��v���pi�o�*���=ϗ&�%�yZ�<I��N�w ���6�\�Z���G�a�����)�$��?���/�M:�
�~���H� c%�hEU�z˛��`�\eռ��B�р��g�X��G�ג��z�ܐ�@���$��=2�o.�@��%φ���(�TQ9z�Qx�d"2��U�saϖ��,��F�2���Y�T�[�yXi�!��=:s��n��{8���O���Y'�4MJh��u"F���n�z�;��w�2\��#{��+�J��D�+m�}/S�J�.]��Z,b	x���m��<x�w`QdjBb�O(��ͧ�S��Aj0��Y��if���V�ڮ�+�K��!�� < ���+��#C�2�C�7����%��dn��N�> y����h�#N��s�mW�2�ɀ�n7���m��;���9��w�c�F��5h3�(=r�k���Q/�qG��l�����������y8lJg��n���A���v�����U2�Y�po���8�JjQRg�������ʾ�fX!��� ��,�u9g� f�l��M5Ln5��{s5� `���5;}z�?YJjp�4ԿG	݃��`��-�.��q#�Ub�_
T�k�S��݄�$OrF��Ata0o!p+�dy�}V��;*�P��&m�z�	i_�������T�{�[��g����in��I{Q����OS�"
n�����z�j�Ӏ�޿���X��(���~X��"�{hM �E��X��yW����[����k����+���Tb�uUģK()J�8�ڜe��k~���Mlz�?�KI�������䔢i�,S%{~[�wѪ�V(�8��|���:����ĸ���
�l��~�2*S�1�\;����`ǅ�ր�ɋ�;ŉ)��tm�6���QT9�T|��W|8ԉ�~?��r�#�Z����C;�M�ꡨ L�;|����Dr[�����7�<灉ҷ�>�� �2�mA�BЕGO�K��;:�b�	x���E�#�H_xVy��-�Jb��P@A`��l��x�"�q�l��9����mxsg��j���CT�7��{��Fy�C����P����/#1�+A_k�=Y�S�a�5���]��r��;�%�����þ�ϖ���mx���(NlPۻ��Ղ�20�+k3�(�l��&�.L�� mD"�C�'W'E���m�_g8��Tf4�����D�M�F`��R$�+�'�a�!����'��=�La6��w�T������r���6������P�<9�U)�smLr����Ӆ����#�����|��s�(��Z�Ĵm��REO ��/�kFO�4���y��u� }�?���pQ��EH�0�b��O���Z6��'�8��O��W/���=��J�~��6I�>?P��Φ(�^�a��C����e��xG�����ڐJ�d��̙��U
�i��g���x���&�=�4���ݝ�D�l��U�Ũ*|���e��;��E��t)�=1l=�X�W�ӭ�6��5�F�
Br��^��G���fv�"�x��ߵ~�Eq)X�[�s��s4���WFs���"/��J���ҁ�9��������MR�
wT�=;a���ﾄ�qm�	�J�r.@��v]�|ݸ�L��S�{%��>�(5^\�dʚ�n��2?�����JD�<��mvoN=�:�<������5��w�W��=Q��rT,�iB�zF�2P'�m���E���f@ w)I����i�gcۘ�w۪�������KA$�\�N`*[�ho�ԾG3IEnS�\�
��AQ�i�J��"m��MM��j�=0Fy�3+7|��Sd;�&#���jb��Y�3FJN�Fܹ9-Ym��pg���-d�yD�D �7����7Z+sEM�8�9L]��C.Wy�� � ��!"^vi_1����cL}�v?�%7{��^ň�R�m�����jC�Ms0D)鳇Z��8
RO�z�ѡG�E�ù��rL'�NX�i-�].�|���/)��ͮ�Y�#���g�♏��XE5^Q�u"�y X����f����)8�@��a�2%k���Q���s8��C����!�:�J�����}Fڦ~z�R��a`1�9	�Pp~��-�5���;����^� o����H�:����(m's�oϲИ%45���Z+/T�)�h ����η>��cCG-��TEKjN#�����&�S�FF2%p��7ԑ3�'I�ac}��!nmܛZd@�vq�"�/��xgۉ�m�� �^zW1��ۛ $QN��|��G�7�ǝ���I���|�b
d���������٫�jqI[Na\@k���g�@���<��#2�~8���v4�ĤR�B�K�0uu0k��)��LT������>x�k��˔����O'�_B�\��~?�M����V�"j�������Ȧ��%E�c������C����s������52���ʶÔ_N���U��aɾ� }�Z���,\���,�h��N��)�^>�I���-�tZa���ނ�|� �)�E欞B��bF�S]QyZ��g%��]	�H�0P�Қ�Z�)����0��SC�GzȊO�ڟtL���S�L���T�W�3q�L?2'��Cp�M�6�]������4ېZ�r!WrX����N����Ng��c���Dr�������fa6�V0~� ���>�ò,;��[�Y�v,�K+�^���`U��*	﹗7�d���WZ���ț�ӟ��Z���B�ȑ� �h�gH���Jd*��2�uEx�u���ƨ����'��c�ٖMOBv��K�ʨ��,�n�J����q���w4�tM�,���l��k�Bg�9c[@c���ىc7���,�
9���|؃$�dwO����q�ǪR����ϟ��/��?�b���������	���G���.�F�g�♰%y��v���+��τ�O�^�):q}�7�����q>��\�A�:J<�gۋ��}�Xu\|5bI3��#�|�������O/3����qK~��o�v���.1�P8&���G����b�J��"GKU���D)�sZ�!*����p�o���X�z#�P޻��&�ىx4����Q�r�`.��0�ʵc�`��B�0�U��sG�<x�xpBVI?���kܡ�G��I��k�.�T�,��9��ӵJ�#󙅬d��.߻�Q����O��n��Xf}�_�}[<��<SD�#K�B��Qu'vp�2Y����`'�l&ʱ�˕I��Ǚ��l��ԍ)�Z۟`C�cL.��B;(gT=�|J���9�;%�X����DnI.%̱,��&%�_�����"�.��"#F�Mq7%��7J�<Sf ���9�9]@8�1X���y��uF!e-�/�c�OW��_َ��@�����I|+�&wGAHj�C������=i�K�E����KGz�{k�ڊ����1aow�������R�v��%��v�*�2�C)����NGv�ޛ� +��V���䋋U3Z�=�U�� �F�Ȍ�W«!