XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ڹ�������ܓޗOE�_�4b]�1��wo+QdCK����*��^�Ҍ�S<a�ǭ�/�ѓuM�`~��aM����ۡ�1�>w����n��):H38�s*�i�'���.�o�y�@=]F�LC_i0��{'G�7��k�͕<�ij�fS�1/�~���(�s�[OR�h΁�&W��nN��I���J�m֊�U��(�b�ْ�V��]-�#�@���k�#>"����Hz��F&�;�}�0�`AJ��1o5풏[�ʶ��"y�cA�~DWT/�&)�(�C&��7-��	�$s�C�n�+2�Ӊk(�y�N�"OFj����lh|��}F��oXQ9e�aG�~���!�y[����j�k'��4n�K�P�P�/=�Q��v)��р�
�,�F[�$"�N��~��i�O�8�� M�Gi����v&��x���u�|�Dѫb���h�������?�ܻ�a��	�ַ��\�lf���wd��1~Ռ����Q�N19Boh"΢�m�N ��?}rj�\��y9\��֞�1M�͟��_�t��^-�&�.hN��!�^ž�3���x��~��}��	1�oP�j��AH��,���M���brd��*��L����ӝSZ!��ӬYPC��!m�(�Oׂ&G��U�/]�8O�ɔ�
�k���S��U��s��w{��B{���RM	2h9/�pL�h�!?Ж��;����1<�|:�#����h�x�(aX#g�k7;:/i��0���R�4ls��+9q�?TPXlxVHYEB    3a46    1050bd��N�����K2��i�UG6�X���5?�1Q��b�}ؠ���$�.�W���s*q{�V��*B�vk���&(${fE��0�Ǹ����?�b�O�5ՌC���?�ܯk�q����d�D1�'��}��s����,ڂ9L<��a�e��]��:�44��\�+����㍀��hl�C0�,�B���
zNX�[>�9T������Ȱ�>l��Cs�,�M�㗥,GW��a��vFi��PH�1��X���qHBU����{����W3�v�ǋ@�2����b��=��C!Z�3ܱ�� +��FZ��9�#X6�-H�,6��c\�SB1R�M snD��emJ	$�{ũ���E�^��|/7�W��� �y0��wzv`z��$˼�+�Zd�}�5A���4W��&� (%��{X���u� ���(�?:xnۥ
��4/t����o�2���ז^i(P�la!9��/�8�������J�i�n?]�.���P@������?��J�fo�����Q���̽S�k�-]�	�2z�����ܲ��ԃ���t0(�K�O�����>�re=lm��k7	'�hz���e��#���bb�I����&O�S$;�21tOܴ�:��+G��}j�t���l�jؐ�Ѩ9��F�Zj�H�[��&51�R�T�i{�I��8��{�2�	�5I�\6�����T��{�,î�^ǁ� ����рV��Z�������ͬ I�`O/В����g~:�J����*�s�d(Hn1�gk0��\V��`g�I���:��y�=w���E�䰒�'�Կ5���aJ��� C1�% �%�����j(TW,f�-���c[s��N��()XxI�w��~S��Q	�l�ۚ��t�������z}y;s��}/��E��ڸs��JH!���I��0+�ֶ���m>�i-CqG=<���.!��� ����o��Ԧp��Y�g@��+X�;OZN�lVv�5m���-H>"��I��A��"�~e���u(��%��L�2?��L4a�62)M�/�P�$#�)j���8 &��ba��0hȓ��r�]�5t�ഋ�˞m�!K��6`�)IA����B�:���-HM�����7h1��G�b<*^�}N����u�_7h�j/bz�h$/bY����c���
�<��#��\�F{=�=�Zډ�����T�MB�E:�"=��F<�L'K觽�C����q��s�ID���[`�ӡ$�P��~1^���h۲.��O[<��/]��E_�{����Q�[��)?�^~�Zq�%�3�����2�a�{�y�Q٢2��c��&��W�)�7q:b���jK�"����V�?�OSÆњ�s��Z���G�շ(\�<��+]�`�� �q�ֿ��$\���`����IOq�?�z[�cVפ4�͘�bE{ ƞ��j�r2gt]�k�w��\�����sÝ�,I��qm~ʸ`r�T�ɂÚrU5g�b�"�bA�u]}趠 Ucm��!�K�n�K}7.��0KTX�D��Ӓk!V�j{4]\V�7�O����ف������{7�h��;\��zէ�_�U����N6�A�{&�v;ņ�x./���۪�Ti�r�x�H�	�`�@o��?��� �6}����z�><��%���Ґ�!�Z�����y���I�)�Oք���򎔨� �u�ۍ{T2�'���aP�j�.T{�1*$�0�s�
<�;��a�Ɠ�:|�߼�������D���M|D؈�J�X-+ ��=�wDZ���,ʰ�!��F�/<�؈�A<6\�@�6[��eC@�ӄ�Y?W��K1S�2��,����s�4IT��<�)L℻�Ö�ޤ���f�7�~S�~*��� p�:BY[Z$��8fV�Nh#�5x�]�j�̏�Y8$ʬ�A��\��Y�#�����2dX���� ��Y#>�����c�*` ��?��r��swV��R�Я����y���W�?��~�x�f1M*�&q\�EI�h�>_�֊�p{�\���_�%;0GeII��E�ez�m��E����b��8��rC��Vu�pm��&y�v	%�8���Lj>M�ܺ�T��e�Y�-�'���_�b��^FK��I���L��������g�8�^�}����|�/W%��.'1�R�jU�enX^���0��S���C�2�ob-	�c��0�k�&��#�9�c:�!�w�S�(�.e�K�H�#R���Ƶŕ�䉝5�&.�Y��HYƌ����O5&$����|��&Ӫ=�b��3�`_z�>�S@�
E��gi&��H��@:14x����hO�⫟����Ka��џkB�Nʦ]|X(�W��_�	�M��#Y3� �}�R�z�����P�����m�~��c&���z-�F��x�2г����/xXm��$띴���X�=���@6�!��W6��u�p�_+�$$z�81p.��&}O8�!F���o%}��b��{��N�ޒ$4$�?L/��&�"a�f��4�(^+�*W**�$����.b}An�@N+�FX/C0<ڞĚ}Z�l-|e�ʈ�'`�ݡ����0�м�)QFW�	)�}�ŭ�}�윤��_�=�@��ـ�T�YT O�C����*?��zl��̚o9,u=�h�M�ճ<��ƙ�e�bn^s�R��sdc��#ރ�[��j�>r��s�r�>D`.�~8hgs�u�V���]�T&Q���B/�Ϣ�*?�g	_{~����>ſ��q��� 骳�;��<��Ij|纫et��Y �h����0T�Af���I��ֆ���cP/�5c�,��AivW_��޶��&Wm%/��U�b5Xu�H���ɾ+-���ETݾ��Oj�W��+�3� ��L�zx��/���b�`Y���h�y�-d�����m�)maY���ބʹ����ecϡ4��t����V�w'������ZbQzz����V�10X4�A9�ZYaZb�~��LSp#�였���S� ��J@��o�,y��E^f�T��4-� ���f-3"@�^���s�,7""��êw��T#�A�M I�I�Y쪬5�E�:a�z�[���/8�{e���`-�w���:�h�(�K�h>AU!#�/ T=��e]�AuMB)�.��e�mS����ZR�\���Z�c�د:������G��H��3GC�AJa�Y����n!a=s����J^���}�&:�)44wK��gV�fD�R��a��v)��KD� ��/�����$	����#�G,۪��?��uB6�*\���3�G,��2:j
l85�4	��7V��>-@��)�cI�N�ݤ��Գ+�����b�!��5Nҿ��sѤ᨟�NU�th��M0Gb���Xw��m�,�4�emQ,fn�@������MVىB�j�t{u`���Y I�[�h�=� ����:�`��Vl_V�d�ŷ��2Y�W%M�\�����a�4�}�N��Bx��cb��7X�Z#�$q^��u���?mǶ1���x_L)�J�N�����c�����(d��2��Vr [�����o&u7聕:��54�π��8N�rS^6�p�EF�=��"����(�Q٬���iV��*lˑ^ǲ��6?RC0���[�������a�Aze��#42��eͦ|'	5�'��"�k�ľ"��s@,�����f�]��,�S�~��I�%�o�J$�Ƃ�K�G0U��\O_;�i�)�;v�T(5���<�P�I����X�:���n�_ S},u�zL�(>GB
1#�i��a' �����:�܄X_�'��V`�KWvsҘy>�B�+c��(jx��$~j�Oz�E 6f�n��k�ۏ7����7�8��򍪰�9 �fְ�*f4��J�l��j��MJ�@0��C� .��K��
N��6���ԍ>|e��>o>����[�����>Y{O�O{���
�2	��_�&[�����nvM���+�
?��ƛ@4�E���K��,��j���J�j�Փ��q���y�a�䚋m��[GEN�t!HF<VT�u�&�-X�ߐU��H�%��J+�ķ�����ֽU$��p�����N=