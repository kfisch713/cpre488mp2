XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n������G��m�y��ٻq4?Ո� 7R�yk˳���g�����=�j&=j��0�v�������m�Mb��:ȷ�#�%�0���b�0x8��E������e�!A�G�T8�Q�S��^6����I�|��^�%�ZLlF�{��6���;�U�������`<�%pS�G�o��~.(�Knn�F�(����~R!#@�vP�6%\��S�Qd��\��x�8-.1�w�6xX��&Kh�O�vV�up$����D�{�d����A�3Py\6�k9�����R�1�s%4l[�*��c�.�/�s4�1�����JTIhZ��Kaj_����T+��������A=��T�P�Ÿ&��ps��k��Jf�00�� �j��O�=���a�dI�|��_�X[8�����/x�6~�+v� �,fWv��[s)�1:��
f���N�K������ Fߺ�}įvHʲ����=��1��R=#�T�U�u�?Z������Z�k=����Z�#"ӻ�~��5FZ�5I��\�[D���S����kǼ	�@��+�\<�����!؊{�d �~�b���j��hwk4�%��'7y�����oM*��]Kn`���I=�L�F��S^��ܷ:��A����F��0���Q�L������9怠7E'<�#s�a���H�q΀�N�t��5zM�+~I�қyy�1{� f����O�y�����c���iY���lԒa���'�)���(�,ԊXlxVHYEB    4284    1110{�������tk�21���\u�х�!r?C��73(,0��cRJ�(�>�=  ��P�����Ԧ��ѐo�aY��Jc��+Ɠ[Z��s1�]��|D�#hs�x<�wT�{�ϡR�� ��lI°<giI�[�.�v�lى�|\��{Y��~ g��&Q�̬��)RDm�8���3�~����[���T�fR]��
1:[�I����Қ��jK��� �HΡr4��Y�:��Z���W5���Y�[��a�b��J���% �w� �?��VI�0�d28���޾Ʃt���x�q��3�VPy�ϰE���HAIU��,�
�Fڊ߾8��<�2.����|���U�^BfD�/�K�����u�2�Sg�gH������MAn�9�>�� �4�;�?������	41��f�qa�'�W�������b�� �Z IͶ$�A2��$ĥ&"_�ܡ�%�>8<���9<��7��h|�6]��R�Q9Ο�%��mw��z�!��e�@v��p*���e����ʾj1�8�����?�;��W�gþiܕ0HS(f��
_Y��v��3�o�6D5u�\4�w!Rjf�|�~kyT�  ���j8����_^�L���d�v�5�\���U���|�dRbE�/�O{mG�U������zң�ᣅ�M, Isȇi�y��W�RK*��������-�~K!�')V�!���ㄫL�Z�Ʈ|�N��J��7�|{��Ȼ��0F_�6�zʞ���c%��{�4�cM�JsG��rI=��;��h[��Rk��K�@��ф�U(l���879����X�(�6z@V�qSe���af�{ ���ϧ��GNU�@���,�9����T¥�eTH����P���&�� B6��Un��펾B*���&g|�j�Y ��Y����-8ϯl��2 �y���ueoF��n8��>��e�7���P3T��X�z;��w6��&z�R�Y�`	P�ېm�n��0g�4^�vW%��L8���Q"���eƥֶ���x�G��98�=�I�?�w��`� ��]�E����2�E��}|��Z�t	�(z��� �e�]�!M��1�n�q���a�k;��0j�^�u��`������ 0Zm�2�|\L,Ce��	n{:�U\;��v��p�r_�
�⿷���H���\;R�rd�&���9���;��d~��������U*������gҎ5�v�Br�D�Qר�,}���fk�3֜)��=Y�O�qJ=�ta�sgFu}%4S���;t�(F�pܑ���r®�ˇ�g�9� s��1Ճ){�O��r%�K� ��}�
K��ɡ	�U0Aؘ�{��v���C);&A7TU��Q�Ho���U�����(�D��-Pg"�ѡ�4���{�k=�Tf��8+�PzϳF�kN}���2z�}ΪYÞW�'C�&�p�����z�;�t�ܿ/[`�ݫ�C�~��$�:��!,��o��c��F�o2��_�����'�e?�e���)8N�.�#��C��9KT����%�k�c�K �Es�ZcsX�0���GZ'����O����`�%)Z�4� ��9�Y̊��%�Q"r�$� �n��9F�H��m�I��I�.[|%�0s��r/���!�A���n�8�xk����y������v�9��G�xR\��)��_������ߐ�ŢYyJ-G˽oA+�kcg��Sc ���^�頟���1�,s&11���jk5���W�3��RVb���a!�MOb]xc5޻�[�}rW�rv	��L��/;�:��Fu���%9K��ZA�j^<��}$;�'ޱ��⧇V�I������7	�Tӫ�[z,�&ICY�� �k�[9�M�bqG��gJ�U�H��/PP"�ր�C2�9���-�xeY����7՜���Sm:"�.�R���|"�l4(V�j3f/U!L/L�e���Tg�Cd"�n����ق�+�s6��Ti�N�w}.c���:o�+L��Kv�)��Q���S��w!��5�67�
��?U��J�#s��Cb�������V��
O�f�rO����
X����8����as$���k]�Ǯ�~OT�5.�g|2.������<�̩?�8ہI'��ص��̿���[.[��A�tN�#RDv}6�֡V~ �,�ᡶ�'��R8�V���X&���L?*a��� '/_�q�M����%P�V������A�*ubr��|F6�o�WLs-������J�����-��&x!S&�� h;h��&��6����&f�+^����� ֥�^�M9�V�<�������*M��@E�m	�S��+�N�Ϧ��4�Ǆ��b��D����<p�*�T^x��bh� �ghN�i�媟�S�QY�ob��U�g�~�%]6#���~U�|]��.��"x�\��dy�>��E����~��F�9��M�B�ٲD�6G�_��p>���k%�a�;Bå�Si���+�.���YWP>uТ)��:��#��4��_`\���n�4|N�逅cF^��z��D�����=�H}^���0���$>�k�x���ª���8��y�JQ�4�����ެ���d�H����Z���6ES��͆��{�|֊�� �"�tXw:`��tw��l;Ktir7�@� +%���~|m�c��^��Q/Zd�����ԍq?B�U��9ڳz������!�_
3=�i�ġ����>�m���ħ �L�S��k*� '(:��$�K�(����?���[������Č�Mo�fN��j]�F�vֶHz�=��U/j���
ыTF:����G�
#d9�qft�Y�9�m�\XVR����b��Di��'n+�^�k$��u< ����t�!�U1b^-a���9qe����8�y�'��
ј��k�b�Q�8#m�k�5��*�ɅaUj+hPaP���-H��!������'�$+�m�<�*1y����4������ʩ<�^������+���c��	f�={NW�wlٚ���?�|��$b�S������L_�.��(I�iki���|J:�L!�D#�ߥKv0�{�"g?��
Xo�2xE��2l7zLQ�|6O�9�N�e{L�6�����/F��b��x��W�W��c���{?]�����GQ���ΈUt�#bT{��'�u߁4�f�B;�)*[���3}��w�'IDT��o�C��\�{�An��v��X� ����$���i22w~$�4IJ�7�;��+���,��:�>�?^jG�@����3���|�%W�̿8�n���n����Ȼ�A��b����[�7�2��萲G$�O*�[baw�+�o��S�>vj��hW�z+�X1�Z3����C��33�B8w�{�m�,.ܭ��(�3���P���`��הz�N���hF�[b�,���A�a6������|�E��{.ʸlH�M�%�Y�?<Qg�8_���H��~�*���e�� QE����|�����{����X	^��)�ۂ*l�Y�U{ŀ��t��y.$Ǵ��Q��@!���B?s^�l��U4���ƍ����Bn�e͗�Cb}������Ӓ�Dv��a�O�J<���]��m�g�<�R���7f�|��������y����� -܃��Ě�jx"��`�L��D��)JJU�dp��(%8�3O�߄y/0��^�VPNU�Co��v���	���c*�Ў�-�mW���,ViZ�:�� �$Wúk�=i)H���r_6x�2U�+���1�mY�4/��l�ǿf!�lɮ�m8��iRha"_vRO�mǭ���J���U8�#�Jk��h>J=�"��=A�c
9hxa �Nk%j)	��G�]�H����^����X�Obu?v4G$��L�.GJ�=�f�-��E�3-O������.��i|lS����)�4$ɯ��W�D۫�j|�bR\���Ӊk��a��x7%�WBQ�;
�$hIG�My�ōX4����*�ب,Vm��_���ig
�Of����6�%�v�V��jּ�_�^���_��!3X��U�����$�z�$c�~\赨��
��U-�~y�i�4k�&���m�T������`�,�0���%�s	�q��X���}��������;��L���*�X���k5�ibFl��ߡ���F�w��߅`� ��pЩ��>���x]�$�^�0��_�Plr;/�FTX4�R�p9�9�P�0yxbFCU=��0��it��(l��$�~��P��$�>c���{����V��{٪�%�AK�