XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J���߻��Ѫ
sQ/Wmz�^/�����C4�*���LS�!]���XF��]#!�22�=6yj\:"��g㹔����h��2����4�P�S�A9�k��oSM�Lo���"On�*r�1�6�+<�Y{��z�g��Џז� ���2���Q����2��'(p�����\\���
�[�f�{Ʒ����H.�*�/6Ч#;⣚q1�o��.x�0��k����K�Q�n���e��W��e���Ү�_��"�Sʫ.f�(�M��Eɻ����8y��8���F���H��T�
4��c�"C�w��)�����ԗ�"Ԭ�W�bt&�.�n�o$V��|΁�?�����������NB�����܀�;�h�K�#���G���O0��ӔO[ؐ ��؆G���_gH�S��kHQ�u����ŷС&���)��Ysb0Hʡ������JH>#3�ɷR���Si��:��� �.Ȯ�P���M����m��r�\Q���%s�AG�B)���B�
!uc#�����1��3TC�@�Z�>�v��`��=vh��ֹt�.L�Y�����o��S�@t#�9:_k#8��:6�����W��NN5D�l����ن�X`���g.g�G`��r,J���!`H��\�&Uŏw+�aqG�E&���������a�g�f����>��PXOɆ]q�5��*��M! �Q] �U& �C�q��{\ɑ�	K�!�S8T)2�"Hoe�� XlxVHYEB    fa00    2040ZN>� nB��0{�KB_,���ɋ͵�>�TA�̢�@�b�'�NqÂ�dP��>{�L�ƙ�g-lگ	w�������;71��{��W���*3aD|���<v�x��:���S 5�1�6�Q�LįP��0��^D��wF�&�K�6�ѻ�R�1(�d�N�s�6�z�t�n%B��Y%���}�U6*ie���X��x�)-o=��i��,9��i�L��T|��R��o���|7{Ԑ��N=3�zB�:[���	���ߊ����yd�_��A�n<�~.��*v��@6��6-	n0AA4�;v6L����y�RW�	�d�ѧMD�RV����)U�$�VZ���{����C�4����(˱�^����1�e�Qy������2�^��$$wq���r�e ��0�m�Ю�&�ԩE���* &k��K��ڏ���o�7�AFП�|�*k�Xl� �
��@�^KԸx���A�ٜ6_��+.����*Ok?��*���-�ϗ/����8�L:�u`�}ɟ��k�aCrhl����n40�s�^vZ��j[|4�H��wЪaK�S	��c�Ǌ�������gj��k��dcჩ��=+���d+�+{D�c~]ƞ���|z�����3���r9�4s��Hc�>I��E���뱥*���YB��"k�)����w�y:b��^�/4�A�ݥ�2y�ROIa�V#�*�J��oTa����3�C0�g�V#5��_�c�GC��>��kB�0�&���Ž���O�Ƹڼ4gVW���<�^����Pr������4�/������*اH�}k��y���لd�y}~W:5�7=Ck��(L��<γ��M��(���	��a.|��
��³4��6vS�A��ѶGǘz�]u�0_ͥ8�
H=��i��\W���MS �� ���:/]��?�s?�Cnv�$e�I,i�����e�ߜe�&
�q����jboO��³|�f�������]��t�=;�Q�7*R��Z�{������~�G	"��JH�G3<j�����/Nya�'���y�J6�=���Jij�k�F�V�4ނ��Y��V]�����mi�&y�kV�~ˉ����U�{�/0Z��n�WQ5���G�O�(�*Q� ����X)&,r�+���+뷉�d#���ӯ�}�<H����hf�E�B�z;�M9�PB|��4���_�XP��1 ��Ͻ��-/E�ݰo���fɁv�O�߼#H�.?�c�Ve��ቪ,�#	#���M =���'�<�������L��=r��k���2�0rB%�����JCw4,�5�s����3�m��Y,�kר6)�(L�P#��s�a����p��ـ����#��G�+��C�����;�L� �p��Vf���G�.f�v��=�&�[���e��&U��	[���k�>zT�X9F���X]:E,�44�ڕ�C5JG֨����EXI߽q0Xxt��#cd3�����ٓ���>d��I$k��?���p�i�u8 ��K�&њ�u<��e7�8`I�Cx�*�ӟ�:y/�o��>e#[%��1��}፲ٷ�xշ���a+�9�-����$�㰴�/#��%N�<>��{���+����git�Ƶ�-�Pa:U��;ӯ�eV5�]��`K��A9͘
�`J�S�x��*
k��KSA�V�0!(�Dcj4��*U��".��K�[NB�u���M@\�}]�F�|��Q��6��/���߿<�ӱ�������B��[/��.Ӻ������UuB��ʫp�f"j�W�4S���:���� ����-U3�V"BGOgЁ�!n�ݐ#�{>Y���Gd$/�<�b�pav�@�g�GB�O]�9��g�H�G2��Xq��;�U����
3��z��#K�%k���5�u$��fegeC���:^��@qo��`4��Dp��a��t�����Ǌ�O╂!;ڔ`P�h�/��h*ݍ�Y����n�r���WSb�� �j�a ~n`:]�Z����-��Ž(0"���ׁ
ߛ��\3ND;�]ڐ<a쑴�&�͕�n�2�Ui֎c�{琔�cz֭�NRƧ� ����O99R��x(5U�,��peRf�����xJ/),�Łd���B�	��(�,��>>�/%�'-�D�P}[�X��v�qN1t��[�n��g%Bs�=qk��"����;"�S�]s�`���9�K�����=o�l���k��$`=�ho���M �6�"o=�R;Q\X��1�z19�DElp�	O���X�e.QŎ����h�ΰS��c�$l�>~w�we�1��|!&�w�\FM��@�S������*�*�H<���"+f�����*���ke�@�?�Gisq��i���a��e�%���=�Th�vP�5��#�z;Pv�Z��G��xx'�����CʸTbA5���%(:��%�����m`�q_=Di���CT��#����������t1t��s&�H���k�]g�8�g!�Ю ��'�$S�<����7&b�<�¤	����!,�{��ŷ�p�ٸ���Fn*d�~s�����kۤ���Z6o�ͺVW��i��Rp��L����e���R�s$������C�0"%z�n��.	?�m��'�ڂu2�R0Ф�L��B:�m T��@"�?Hc8�(�P��|�ӌ����zZC����*�h�Yu��4��T��=p�9�F�D�L�%�q�n9�S�b�5d��~96�mup�C�uY������1�c����vi��������������bY#���[�A�x���v���V"ʙ� �Wٙ����,Ŵas�q���� Q5�X�LȲ~������e5��!�8ގ���ң)I��֛��BZ<����V��)�(��#����x�bV���d��q��Eԛ�WJ;�_��5_x��B �a��?v���Oo����P�;�k�[�����,��QV�L�E��j*J�tHZ�k�jv�c�X��j=)U,�٬D7fp ��*��t�d�\��;��(^�
@04T�.�u3��E���A���$1�؈� �)���E�ά����O/>�t���Q����+�ә��� �ɚuJ�= 	�_�b�
gG��`�P'��n!XT��
��~ɇ��,0Ӽ ��Nԧ0�y�#pff�b6B�2�N�[^M�ҩOo���'�˓��G%��?OM�[#ˌUW�T�
�S�ܬ}1Z�d!+��z{��K�a�� dc��Hd�)�K�3�L����$t�R���E
@ZՉ��kcΣ�o�jy"D[VZ;��i�B��S��~?��3�VV¹߽����f�_rk�I�D%2�KW��mx>[�jǋ��xT��@��B��/���h?�|8����8<�͕H����Vނ�<J1;�c�[�&�����UU�O��6con����bwD��) _���J��Ž7�3'!�����^���ؒ+�v��n�1{��cG3��[t�"��f��ғh�L��G�S;p��d�����?��`"�a$A�8�e\�e_��4���ew���X왽�t�Xh3�EL/O�:fV����ӌ�hOe6t�.Kޕ�
���-0�~Y%��+�HT����E2��)�eR tL�u�# ���p�r�&3�A��3���B��]=��ls'��I���ѕf8�v"�mV�3��{�$A�r���~��	��H"� (Z7%��":��ܛ�������N_U�s�{V�&ֿ��5��bR?ٛ2�࿅����lq�.��&���u�W��R��=`X��բy�o�r{��Ҝ�TL'2�
�j���BPdhÅ��Ș�;��(��\��H&�)�7��O|�]4��b����]�WB�)(؆R�	Ny�N���Mw�!!]�-��m��`�W�X�{a~��zYC�	�yܡ.��h���Дo�*��R��4�	��b�h�V��+W�}f1�1҆�>�ၝ	�����?���mC+��m������h��Q��l���O��sg�Ni2Qx�F�f�fd�d�Mj��ܤ	�Nr}��L�UF�!��A�&�ɷ�5��1-j}W���1�"6U��ۿ���6=���0��[Y�fi��?MD��5}���!2!"�+Y.?����<edsmD�M���t�m�qA~D��2[�Ẳ��0�eQ��������=���6��İ��� ����A�d���o�a�PRF|�R�O��%�K�����z����?�Y,��"�ʆ<V<���P~�Ec��|��*k�g�/
4�H�MvKM�rTQ�z9&�j2��|@)���A���=��r&��]k7��C�%z�����3��`܏�MT�o�}�K{�\��h6Ӹ�u����L��X詉��!O��e�h3��q`2Oe}J�Jְ*��G��e`���"���D�p�Þ�^xN�$��+ ����nY����t�f��ޝ]�vC_c�?���b��RҦͱO�?U�@�>��}"��u�lAN��9��?�/ޒ�_��4����i�!�*
>19e�� �&�����4�YuW� �]�x�Oژ+��󖎉-	�k�Ȼ����O�U�$t�_��3���;LXYkSP�$�L�����yJ9��̊�u}º���v�GLQ�:�h1��K�`���O���/�ƅn�z�L��.�[S{!;�����G�� 9��n�".�g[8|y��[9�D)=�v�:N�k�:Pq$T��@�4*�P�V*�0��R�@k:�˟_���3��gH���2v �;�~ſ$ȷ;��/e��We�Ŗ���w~�A������9� _d�wJ��l?���duui�nDc���$���AL.�f�lO����abEUa�$#:�봈1O&��4O�%�EW�߿!�,Q��{ej��\-����,"�L�@�L��bU���"k{�3G՜x,S9
�i#��7�<Ut�݆���(���w�T�_��-.2�}���ϔS}����-~�$�{DE!�O��c��ߠ�7,0��d�Ӏ��uy���1g�D|�D���r$��y'�[p�*c�l�?Y�<����d�z�T��[d�#�v�>{ӎ��>Iئb���s!�X�Ar�ַ� ��C���^�Ip��ƚ�a5?�������~z���M������g�q1ڀ��䘬_g�9mt�`o���2-��B�g�cdt�oZ�ܧ���g�.�)P];:�ڤ���,xCy%{��_���%�=�X�c	W�R��d��+�R�
i	^����WP̿����jF�'���P!�4	x����{s'a��;�G&S�g�e�1�W:�kil!�#}ߠ��^�M��U2���X�sh�;"p~�QW�]|�,C�ޘv�I�lvTNv�����J�F2p��r��PU�dt�p�ƿ5YR�Bs\4��B�.9�u�JrM�ZͼI������ �|\�W�K
q�9;�:��n|���˕�Q��w���Y��<��-4e&�4�Y\B-�!tb��9]]Z+�o�E�dx�> 2���q�<=6�X�J����a��	T��oדUb�}���͋@:sS�g�\\+�C���2�3@#v\�ݪg���P ��q2����Ь�J4g�Ɔ�Ȣj�=����B���H���C�%ug�E>{�*8�O�w"���]�ubo�7 6��1.��;Q�;\��Q%����c�ٺ�9��~�=c�D)�SƋbQg��1;5���3
�4��ۘn��}N_����}���-�o-u��"�ղ�"����P�L���?��g���H���<l�_k��S�Ƴ��^�hz��]�7�z��y-�^��v(g=P�M�����Yi�o��ճ�V���?m���>��QS
z��}B�wu� ���r���I��^(*G�e�y4��qo������>�x��=��otKT
[�S撆喠�D��l&v0�7C�eO�ĝ~t����5E��K�9!OR�ƒ���FUTO���]�^}ѩy�G�ӯ�BK�a�uM����䚚�q�'��lt���Z:��E�����������4�iƷB!�݂�G�[tm��;��X��w�j\��4���&�����y���Z��l�;U!E�@2M�e9ئ +�3;��Y��;�PE��MV���+4$=�Z����o���.(�%SU�Ot�(�CV�F��vWz!�dG�.V��w�WUQ��<"���7w��N֩��5@����	�r��ڽ��}΂��mę��%h�7j�r���q���(����.@���f5�u�_ K��z;Xȧ^�J��H��ͺ�`� *���-��Ǥq^�4��p��@����e���\nQ���
\�z�f��+��y�C��#ԓw>�i �g�&����n�<���e��3�^����d�.2�㬝�b�q��5�
��P���p� �uR�@�L���eٌ�4�}N���h9�������*M
t"c�������h�2�����?:P��&z���!��N`�XxtAϜwJ<[�50��v�L�\��4y0���[s���M�(Z��+.rt��A����ڠ{�wG��Bk�T0���9l
&�}�6���`##��_�z:�#�
;|,SJ�j��S*$���/�����.���l�|#�}r� *G����r�W(T��%��3d���v!x��kB�Pw��������L\T�_k#�����w�rڼ�w�����t����W�<_�1�k.s���e�viEo~�!�@jX�<��ܻ�GS�����N.s��@T;���듪h�[ ��h�X�$i&@۹� c�ׄ=}_S50��x�=G4'.2�rv�����+�v����v��Z�T�u�q={t���^Ͳ^���vh����ѫ���*^>vr]Zw��f%ؘ����ٚ���
��D(%�}T��N�pT���\�� �LQ��"���A}.X��o/�[ma�"��G��1��W��~���%�0�u�5F�B�9�9���{>��ʚ���s�7r߸[��֚���q��d�j��tGήBZ��ӆL����$�����bB���})�3ce����x��]�����gcL ��D����I������gpd��)R1|���+�U.�J��3�����b��z>8/Ŧ��Ĉ��i8i���L����U@��[�϶�x�}��7nc��{sGs�����޹ �0������TOT�S���@0EB����Y}�s�w�����(�#���f��/Ʈ%L�6l�ii����B����"����+,��4�G(�fa Θë�����]�e���uZH�X;W��ɕ �y���!����-+%D�Z�#/(���4$,REV�я�����c"TժK@\/ ������"��4�g��8����.6_���E�GŎ���d�&�l磊6q�*y��=e.���Q��}�������<b�����D�>Pc���b�9V�_�a
���h�6��`3yW<�KΕz������~�	Hn��@{N'$��(+��^��
�sj�6�A��*�ë���[ �gyv�ff��Y��'��(��	���	����sՄ�	;H�1��x��)p�$���*�i�+x�(�4��K�Ge[">-@���q%Mj���t�qE@T���M������\笤�㙫7�%��
thV��}�
N.����d@T�v|cq�f$�j��0��m�5��� �T\�8�Z���+*��?�?d�wv���)XTnZ;E�.|8��R9b�1���m���ᆸ����3�<F*Zd?a�h^F�Lt������+�pۋ��I�	_�.��4��I�<�"ٛ�	p�A��&g�aj���r���o�v�__w���D������ej�b�e��g}�x��ퟢ�$A;_���ˊS��MڃRR��
r��8U�g�s��+%9[br(D�B{n7���K �",���� +�2f��S}�J�ƴ	���Z��!�+�o����ne�'3�7�K��h��$������:�m�n��UFjԩ/\�Bﰦoa�:�-l��q`$�
������M5�r@���sd�}��4�n���:<�t~�|��a������@;�aد�9R&V5~`#n��)*xN����Pߙ� AѹWf�HXlxVHYEB    4f62     b50��dl�{)c��@�G|�ĦS"��Z��J�^BHoD��UaC��)W�Hz~wC��\a��0�&T��J�D3����5o��B̎M�^�]������'���i��%�c�q$:��_S�ρ*wˤTǋ'!��UͲ3e�E���P�v�~o�����8�vHH�>&���s�`;@ܢ�3�eצf�%��cDmo���@ߠqf�;�g�*�����0_H�3�cX�Z�s�Z�Uy<�]�6��c�^���������@�W��ْ���7�_�q�ol^����q{PB����0 �xc�.f���3:$�K﷧�`#Ie�8� ��̽](��VLVY�"Ϥy�ZX`�N�]��:?����5w� `����!���&VN)V � *>(�=XHY\�:�����h��-#}A9�(��	���J��imMN1��df�EMnު�k��54��[$.e�/��]!�������={ Q�*�Т6��O.|L,P�F��I]�¨	h��u_�JW9� ��Hu�ޝ�Vb9.N�R�Ca�����g��7��I~��z��"�c�*�h���'0HÆ�A�"�ëo��ͪ�KE��f���`�X��x�Ո�	��r�6�AX���zԳ��we�m����x;���ݢ�|\�yF<������6���e$��)�W	�Y�,}>f�.΄FQ]u�.QA��l��Gȭ��Y�*8�n�j_Y �I"�y�cIA��+����I�%�rF�����}�j���4��B�;?�&�F@k�a˔(m���av�|Ε��x�����>�O��:�f���,@#���n"lA�-"�'`	�m��2vD�Ecn��=i�v��&�t�q��-b���9q[�JU"�,XR)��7^�u�3Ģ2@���A3�7'��YWl<�|"9�B��l��2�'��h�<^�+��=_�9��d��s�N+�<�*��LlA��	.�cu�F*�f���YG�&5 Hd�<W1]��Fb`��0-壂	���O#�e nS�s�(�dhn�Jo=,3&f9�����A+�^}�ӊ�/�@�"K�*A՗�X}��X��^�xKw��I5��$��Ɂ/(ؠID�~��PU�'lO�Ybv$�����Cي�,$�>�9�J#tIEXZu�T�:�8	m�(��0Ӗ��(��Y�{���vPh.��t�#��dݹ���.Q�=���H;�����A!�bf$w$i��nL�5�� U?Ҩ�v�>;ަ�E�� ���f@�������q�f_�� ��?x�K^�(2�u�N��f]��gy����0� `�������2�#u)�%�͊h�J���¿�����z��UE̽u Y�ZY��XZ)�eI���{�@W7�֨�N���P
T)g�,h�R���kHIO�ϤTL,O��ǖ�����EC ��w��K� q1���g���94���T��x}.ΑF[7���p��(
�:}Mx_!ʱy���=E�"�>�*�ݕ�=�� �z��/Ӽ�ؑV��%��A/ª��mkh�ٖp�eE��B9�{�*��8skȎ��!	�>��*z�{x%�xW�`u���bR��ͽi���Ζ��k���"[�@�����1g§�n�B������Î(>�]�%%r�R��g͐!n�b���J�D�{�ggʹB���Yc��;�Ai=��7�v?R�w�Bʞyk�XE;�LEZbU��(܀��p��6D���:�W��d?�D"+�."�k�R��3%S������s��Ζ�<�O���n\k�e�,`J/��	�M@H،�+[_Ik3��'דn��>ޘ�b�b��X�ڂQ=����<_4�x\l�㗠�`iL�Y���ZR]x�HN����WE��wӗXV�dt�)�V����u���{:j�eh$�AC�3b��j�.>,�,"���n0k�ZOV}?h�F�U[=���4�8��>A�-���}���Y!��R�LW�U�_*�h��!�S��wn;���u��%�����;Uop�1���l�6�K�'|�[����)J���C��	�d��'�`�C��L� ��4�x��_����J�g �h�2 �Ǹ��W�F��6��	h�Gl}��y���K+��4t�Jf4An�͑��c�I�pA����J�F3�:Ov�>.��J�%FqSsB$��۰��t��	��������U:3ϛHѺ$��Է�������Wݷ��M�0�Y�㨩�JJyt�/����4�P�j_�:>6`nLw�)��T����\�ߡ`M��S��3��Φ�1��Gp�Yě�{Kޑ���1c�������Jqy}�7�;�����e��;������@0��e^b����7-�#�S�q�}Ad��^��Q+�� 6[�oI�n��+�q��e*���ￓm
���G��e|���!R����͜�AR<_sF��@�Rz��e�ˋ�%O�����G�{�N�yK��C4���~W���̩9��vŮB���2Z�H�s�q��.�2@�.���Ze�U}Q	�� �~�=��6���[���K��p��Po�O�yR<Y�R��ɢ. ��yS��`��o&�Y���6Q�b��fljѳ���3�*e�bX0AHw �}S^�������q���M��)K����wڳs �b�d��Ò���8hGW�5�z���x�?�Eª�_���r�DOt��մb���v��C�B �r��������;�5K��,���x~K%����#�G��U[ԦF�07u���0SR7��"Yt��z�Z�-�0#�ɞ� L�cW��#��Vj�4�p۔4�NH[�� ��8��btn:���.!ͯŞbr�ehE����h�nV�� X,�j"�㍛��ٽ7��f-m��:ۈW+b�#�[�x����\�O