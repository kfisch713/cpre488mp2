XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'/���RvO�\ ��_���^��R3Ʀ��?~#�E4[�*fE�ۺ�x5�h[j��,�u��<;���<G>�N�R��{6���{��{up��}5��x�s<�#��-��Y�r�XՑ��_��F�� ����ג�T��P�*�%q1�'{ ;�9��kpԳh��.7�q����(�N,�r����9� ���;K��60Fܲ���R16��j3,��˩j7J1��|y���.=Sf���I�y&l,��EWdx��vf~�wü����L�N��`��~D׍�(.�*��B� �bE��Z���	�>$/F���ξ���A���U�eM���?�y�H��ä�	���^�0y�886j�'��.l4j���,���Ӏ>h����i @�R�I~Y'��A�Qn^F|`��NӶ�?U��Fe�,0M=�ޘU"�'8ͱ�4z^�p��� g1RM�uD��XY�K�q�ÉM�%��C'��l!� �Q�hd�����13>0�"�!�-��9w�������,ȇ�4���B�qcWB�BO��j%��wY�L�}��aSg��
�)�b��Y1y�<Ϸ��v�L`(:]��?4�^����ػ����mm�� }�k��Ė�\%W��8��xI�O
�F׆�tL���G!�p>����ŕTG4o:F�=Sc�Wp��/��1F�^��#�)H�V���<�&�h�tT �D�4�&t?��x�5��g��#�Z�=��J}�~��і�pa\�c/)�)�&�(XlxVHYEB     e07     680�������
�hE9���O��,�W��hi��A
�ݘeWqlU���{ۘl�E�6������J�YңA�g�M؝6hG(kij��<�r'��@�~��ā;��[�]$����n@���UC�H�6��K�	Oa.��>��H��0���⦨H���^���o��}V�f�Y�^�2�򎞱��7x���PN{o��sc�5M������N����Z�g3`p�)�ys�Oo/Lv���C�GL��ez���bH�F��n�jK�l�ʸ"�2;�>��_�3ֶɍO�B�2��̏C�n�~;��a1?D>>\ �v�
��n�r�ª��'��(f˺��I0಴�*���?$o���n��i���b��$�Ц����
�>�i��֧h�� �Y��p��˅ۍh�	�@��U�l����� GF-i��>k>��]��<!?uYڳF� �o".2A�)���-e�x~� �0��	s�I߈���p���y�ս9�vV�wZ�i䦐n2��ipd�Mw���� �ǀ���wd�����nG���Y����!_[��j2�j-��ꭅmg1%Wze1`��\]��R�D��������	g���g��jx�狴�b�ܭr�'�@�$��������Fd%fl��@�߿�@�r'#?l)��	A�.�7L�����	�GǕ ����w���ٮ��гZ�ҫ�ܐ�W{,��g�z<8����L9�%|)��e��LN,f^j�{ґ�������8�*��"Z����hދ���M�����áU�I
2���~2�k������}����Lڤ��B]hS�H��L%AP��^c)���YN�8I�^����!�S�PlH��h$��;�S��M�M-K��S��ؔ�sQ(L�ro�}5*0~M
�h��(ւ1��I��
-	��ʐJ5BM%�^3���t�K �[r=X�p�<A�ɳ8�ƫ��>Iil��-�ܪ@F�$��#�<�X����r��갽��;}��}U�>0d}�\	�=��J��@�)'m2��0L�)>.7��ky]�V��c��뽮n���&Ӆ=D{��QQ������cq7$�s�}����@0�
�z%sL�$\Cw�W�ͅ���M%8�&���4�����yB�o�W�Z��};6�/:[[��n��=%�=WK�ҩy��GV�;�C�rr��yvR�_�2�U%+w�.�Y��	���a$QH�⩫�]խ�V����'���F�^F��?p�`ukM�$KOMR�)Ƿ�:�I�(�O"���Ȕ��č(�M�4=�,�$�z �o�	�0�o6�+;�"4p8���q��%�c��!���2Ec�-S�afA  �ӕ����d����,����aj����OӐl,"zAe]��<�t�W�y)%J������W����+�8P��*��E�w��P�mEX!���B�)���gI"��L�$�GGɲARZ#�}�ËR��Y��ݓ���u�Dj���vk�z���0=Q}�*|�?q�'���7�J�&���2,��]:���o��/&�$�����z���k�;�_�s�BK�������		0�!F��U��,�I�i�\��b=6M�%J�;?���