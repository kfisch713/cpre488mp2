XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����@����6����]sU�� vnڹ6A��;�=�$�U�r�2�S\l�����y=��F�uG�p8��Z<{$��];�:�%_Vb��c�"����G�*z/&��c+B��Xwl�.:���}ʣ�k(�D�w���i`;�N���8�nǻ� bL��RoC�]fpq5\���h�1d���p|����Z}�kƍ\�fXo!Qu�����)p�w��^
L1C�󼅉���<+r���:c��r���OS��sJd�b""=���gf���K/�
Y�?x�i�rz��j�����k"����?4@HǦ��F_G�|S��Z����\���w���a���Ail�م=?��6��y�yYōxZ�m���9�b�����W��m�3�j�:R�3��܏���n��i� p��;�����:�_<`5v��7�o?M�'j\������ �BF��i�7�{�KG�Kr �;C��K����+���+��)`�u�ݡ>|a��f}6݂
��̯�5���ݹ�r�c�� y�Tu7��5$Dz����� :��ڜn���6ޯ^�+����a"
�`����s��b��{\�ފ��!
��D����ȁԚ��Ԝ����@p�ڨ�j�Lټ��]�삝1�GP8$8#0ػ��L�\��m=ꓪЍ�������z�M�ט"���U���IL��\G�Ͱ.��8?+����l?Y&��*Ć��ջ\QW�1����^z�%�G���oXlxVHYEB    1a34     990�f��B*,�Fon��diE���on�����א��Y����������\��ʶ��=�XJ�Ծ�`6y�iW3�!U�q���Ő�i�[ n��Գe��*a���?�w�f񐪡6�n�I�O��"{Ay5�k�IC�['�S�VY#W��d�6Do���sR�T���]�^f���S�EQ�s�ON#P�PG|@�%�� \˶8�;j� �>�}�﹵�~Vy_�⫝̸����h
g�[xC���"em��l��(:�89��iy �nɻ�Qͯ�>�(m�n��yx���?$Fj���/c��N�:P�u-�]Z�F�@��0(��'!>L'�ڹ�}�YBbU����-���d��o"�7�,���n��?(�_ �\n��h�6�'��BeOF�~�J���K�6� .YӍ?���"��)����7S�|$�q�x��	���y�t���8�2��7Nĉ�6�}��a��)��I��!��q���t��l��"j߶��>��=�I<:�ʋ��̋h�$d� A j�o0ZfT�Մ�z�{�:�5_cvu�p3 �#��pyB�����_�D؜i�q��`(F0�%��PV�� R�"�xjV���b�`�7����l,��1��Q�p��d�9�T�f^�m���1c����fԄ�a�l�X����x�_x��<�mQ�u��&����ؘ�6K7�,GC\���3k�i���)��=V8��6!���qG)[�G��m����R��H��-���$S�0d�s38x���9d[՜�e������r�)��~1!o3���}d�m肓7c�V�͕t��kISE�|ޅ�h�K8�T�~lzu�*H^��<l~��C�B�1�*�.�����8r\<!� | �z�v��rI+�=�,�82P �_vՂJ"�J�+l��w�)�$�|���Oil�<��$X�T0~	��a�jH>��3�p,PO��ܣm_�NB����K_�TYK�	1	����w��w@߃mv�;�y�(Ŏ��� �h�V���axU�l��=W�=�09�3Se�X��o�^�����T�G�c�2�����I�߆�qgǓ}��C?K���?h�#OWH�jU�#��}Wֿ�p�)֙�$��0dcN׏�@��Q+�<��'�k�aO�Y�Ԫ�p_�2Uf>��x�ך%����j3�"�}��[h��u��覢(Hu#p:;C�~e��ei�^����*lb�%y�������EQ������՝���NKk�Sq�*��}��\vV7�!&�l�v/8?d"�3�P�W7��Z&�E�����<��!{%���u�����<�F'�>f�Ӷvd���$\��@XF��|�w���~t�G╒WGj��\u���\,{*�U�����m]�Ky7RL<6l�����O�)	��ZI�YsT$�}��4L7�6[}C��Z�����C#vX��8�����TO�1.crj_������^/�Z��\_`�]/p���p���C;(�1=)�J�9�x�9O�S&!�Țh5\2GP�aat�m��F�v��c�3&�?$,%�H���%\�S��VQU]M����eM����%�qVA.��v'ΑJ`�]�☳��r�ٹ�ⷷS�n�g��d�-ivR�����ׅ���fbG�Lǋ�9{l�`E�1ZqN�A�)4�Nnٺ�H���ro��M�J�<���x�u)�ai�g���.���.m3J�d3����_�О£g��G
���m��y�\��6ұ�#�<���!6��I�
b�Ɗ���H1UUG<�s�U�=��GR!���1^�s-���K�
�����XS�NS�')�򴻽WG��2ZH���o/�����L��:�w��#<!V�с��臱�v�@a� �D�)8���T��4�ZmBXw[s�9�� �Ef��j�]��r�mHVP�͓�3_���@����љ�$�+C_��黜���_G�T��{eU�)�&?�_D1]�,��v���c��5rۛf����_��~W���×��tv�GMwr������i����Я?H�J��G
��Hw,A�	�d�k# U��Ǎ�@���B�kr���M�Y?��P�~��x�x�>5��¥�xx`P0���$'�����٬}D8�Ef��І��F�[�Rؚ�����js�鏵�{�h
��Q9����Ȳ�m-Ml��� �ݔk)>��2������XcaWO��,lp©E��53b��}�)5g��φ�˥�u���S{"8p�-�@h�h�d 	zLk� �{���FC�����M�q/���J�����l�����)O]��"?�#�=�ADK);�A�*RN�&T�D�0*̔D�}8�&2\d�*��I�b�vKVba��M�X�pO>W��L�:�����~�ۓ�f��ϼNO��0ͥ� ��c ��J?�WGCFDB^��'