XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���w�L:���%�g��#�����cL7(��+(��Y��?@�L���?	�~�	s���2���R~����77�CF�o��x���`�d����N�xŮ\qෝ:��*�����)\��ͮ�G-������MO�*L�,�j���Ny��^��2
��;e�I�K����?e��"��E<!NO��r���'$��w�_��WJ�q��-�����۩�S��m�� G~�Q��{v�?�g#�Z�s�����~����.�&���y�w�7eǈ�گ�ڒ�gB�'&ǵ����)/�b���D�7*��s�@Bw���|\:�(��XТ���*�O��3������5U�Jry����}:[i���I�]��� �i�yי��	�������?Ԍ����M<
k��Ԓ@�%Q��,x��;��>^��`���=]�>��:*�Q꾲 �`�h����;c�=f�IQ@�"��f��2:-q�/K��0��׹���l��w�0�yV�f�>gː�A����"��Mfn&�)pf�cj<��H���l�'k��~'[�9�3���Zm�qK�hJ�pi^�'��3�OZ��^�V�Ҫ��������yixF��-@'`��,"����~����?��:�V�Ӑ,�lH= ���x*��棪�i�I� 
=��F��x�.;0��A����;��V�a'`���O<���K�7���Vg���F�T���M+��x�Zֻ,.��XlxVHYEB    925c    1a60��Ħ���)�'L8$�c��%��8�#^�g8%��N
PR-�W���i��P�ǒ�=���f����rg�����]��|:�V/������~�;oIj�V�ց`R`��'X�[���G;/K<ވ*�s-�	G������)8(��E���A�κ�g3���]��E�o�qM��%��V�������)���C;꾩3�zk�?0K�5�S��
~)���Z�;#���=٭����\7C��� �8::N;�$&����a�l�zG��B�6&^�fEo�Op�ծ֗�� ����^ts ~Td|�w��L��E�D�5Z5�x�U���
p0��|�&��	�DҜF�7陴�O n�V1�)y?��~��������P��yaHZ��#&�������FA:�gaX�.kf���+
�i	Nu�3�
��������qr�lK�	�~�@�����C�F�B���O^I��Fw���Z�]h�T܍% t#�@H�1�3MI��K���mo��� %iOeJ('Wor16�K��ۮ�qo<���eU�:	st��*s��cEܚ�����'��Y5��E��a^���i��/�db��/I,4 �i	�0��&�2�������(f���zy�Fk�A�	�4� }��z�WVW�ُD<o��>sT)�5�f&0?�WϺ���3=� �HJbR��~�p��RA���s��!�?"�%�\��m�	�����VZU��N� I��p}��wJ�cE��N�{qƑ�����;�I�V�Hj�!y���#�Q�Ł��R�i�r��]M!�;1����-��y����A!�g���ɝt��=&��3-�%F�wLY2�<d*���u��}�#U}N�#6�[��}�	Y��$Ț�&�_��i,,�:
6@%�#h������>샐�s�X�2�U��I-��j:Ê���U#�9�ګ�Ց��x"��-x�q��I�)���P�^���ZV������b߮6����iqL��k��Y=����ƪ ��cZ��N�H��ڬ}�"��J�Y3]L�aX\�a���$Bz� "�!?���_�Yo��.�+2
;*T��Y��:,$�vg�Oo�����N�\��c�!�I�쾰-E�m�m�i��c��m��5�,���]�!]���"u@��Q�}��zJ�}"�TQH1P�}�F��0^�p[R�e��m��W�Wyya�<�}���TV,2�bc:m-�����;.���[qϭ�dx^=3�MrT62�={���<Ⱦ�gCVcS��dFP����K{_,H�O.^���ǖ�s�~��t���Pf���h�J��K�Z4��v	�������`�;��ix��|�J�y%��^�O@�2��i�xj������ӆMz��cgk�|k�h�g,# ���[�h)��|Y$��h��p��2����B��>F��T1�A�J;�j�*s��yv�;VT�ls�Uc��^��^?��=��y}�R�Hx���$Mw5�8��1�N�73�C���B��,��Y�<��gj:�{�J��_PHJ������7^[��U�z�ݮ6=Τ*�e��]�����;���BzS���^)>P��9D��d�R`�ł`F�sG���tI����F;v�ؐ��c�M�2X��s�:�,z�������{u�}�s ���Co,�5���uu!/�� +p�����cZ���J\�t�/�0�����lB��ƞ�1���{�n4C���)
�L$���a�¥��ߑg�F����䑋i�����R�Ϣ�Ύ��B=ڟE��� �b!@R���ѽ��S�!��b�Dr�KB��E0�.+��Q��0�����=�G�Ͷn/.@��2�T.�{	v�q���8&
���/�
��N� 1:��Q,�|���B���w
-�m����
��V��O �����9�M�̤e���HϢ]*��d��T�dMQ<[}��ɢ���4��@���W{?�s����Y)�lk<�L�4BH��S�X�j��|Q��'�m��M���$��Y���u�.*l����{肏lTo�_߂�A
X��/|�X�m_~� =�ĺׯ�PF�2��EA�t���2ڛ�%o4��#/M�ܖ*��׷����(�KFpVG<�ő(r��> +�M�&�}�=�o��|\D�(RFf'Z#���˄ܔ��^��r拣1vL���R`�T�elln�L��?�_�h<����>�j��?_S�!��Cn˓ధȄ>������tDv_�ଝo��� 8(���Z���T��F`��-D\+CM������I��֐#.�'�.a��M�8�4�l��'ڨ*��(����� O��1��gEix�-�$�f�g� ��v�豑�F�T�A</�,2*���bjm������b�=�x E�[�n�~ �õx����s6K؜����}279���s��tY[˦���L�(M��5�5��9��h:���Vɐ�����<��t�[+#�^��i-)���1�?��ҍ9�E��w^�Uԃ�����([ȫ�O������=����@��U���nY	��)�(���[a�rq��67���G�x~���~���d�E3K�N�HD=�7m��|x)��6�'Q\N���ʀ]�I�)!��`B����U���{d8�}�Pv=�]j���@v�d�
���;�q6 %�'GL��Q��b.�	@a�i���	�_
 �~�ٲ[z�UJN�j^y��=r�/�Զ���?DK���v[�m�p3�U0��j�U�h��1F+'�6& �H]x��=��*)}/le_]=S�_7�-��!N��e:";}c+#�����OB��֦��r���P���_Դ�!��u�aB�}�qE�ſD(�?�
�!m"O��,"4���GҖ�Q�������jb#���y���c�;k�7�n�g͌X@�����O�M�ᕊΣA���f� �����bD��`�~��l�o:����T�VDS?e�K�Ybzc��B+�]8��~!̀�Bh�>0��WYI���]�;��~��"��yWB��x�p���H������DB�b�\g�^� �9��|�a��xp�
��3ǌ�*@+���s�/�!�6T�˔h�`��žk�8��h�S�Cw�����u8�wEg6-x���Oo�c_��(�oa�̻�~W���$3:f�m'�rZ�_�T�q�LUn*l�e葑����2�(
��r�T�B�"[�D���@�l��b.��:�%�1�_���l�I��o^J�"GA|��������S{�C�1�����QO�t���q�\m#�jUE;��h��B����0�J'�
[?��J��P�] �i�Q������'L�^��&��(�f#9�_��+Dr&G4z�Y�Jv���7��,��k���1��F%��;��(�J3�(oΖ7�����A4�&S��G���:<�_E��[QV����"���T�B*Q`N��Q��@Mg}�b�7�d�Ȫ�҉[�Xw�.M���{߹�m�	���a���a �c�sS$���r��=��6�\8~��u/k�|�m��<��`b�!Ŋ�[QŶ�N�?Q�F`R	���~޳f����&�͐���\3�(�^7��D�Kq�g���C-e:L/����}�h�1����1{kJj�k��ɉ����J__k�P��1�ݰI�檸�霸ӥ��6�+Db�5	�/Q�	�x�Ŭ����	bg�� Ҋ�ig����O:��:�L��#�dUr�U�c���
獙�8kl8�S�I�͵�0n}�hr��O~�j�i���C�䱸�3ҫ,�}���Ӹ00.��.��ב�* ��.K��sU�P����q��9����x�GZ�����k�y>f��Y�~�'Tjӛw�Wh�d@�[{x��e������{{&�l�Vj_��3�6�+Z�W��FB��9O]2ꄋ�h��K��0z]�JG3�K�������
2�W�
4RE����[\�-�v�A���ɟzvb�-b��� �<�~3�7�B"��I0W@*�k��Hf��!H�'�$t�}�Tv�qX]�#Ո'V���D鐓O#&�L�4:I���9�.Y�VQ�OX�^䠿�q+ɝZ#)x�-�)_������+~L�p��+ �a�HvMqN4�;]����%/Y��m�7��vƾ��c�^7������ 6.`?%�bU!���n�{�� ����2-�q�a��%�V�d�4�-���<cT�̑=sDP.R�n�Z�*DӬ�f,�DY񋀷�H�02"��-�3/�(Ij4���/C�%�<�l"��qA$g��%������i$� ��-��+��%P��2Z ׭� 8��ڍ�FKnF�Ui���G"�?2�q����/G���dܣB��<R�Ͳ>�ȥ���2'ܖ�P�Q@�i�!�+!�ft��c�0��	�om��1����6�}T5=)a���6��l��������97��E/�zZ�8,���,Ivd}���c�W�Ór�vD|X��l��6���ӑM�"BLb�=�	~�Ba5|�a���5cuGBH.t�!�I�:��I�l6��v��H0�Pm��E$AA0Ą[iacj?a�B^�ޠ2"�HҦ�Mc�)uUO�)]�DΝ��!?V��?���"��&�'G�}8᜺:�ϴ���.�Ե�O��_�E(?��Ƶd���k���R�R�@M
�%۸��Yp���� 9 ��߫�#ʶ�.����4J�����
�o���t�>yz��cq���������tD��2w����i|�,������֩5��wZ����y[~d�\�C��� ��ǹ��78�y<X�p�o���W��MV#&[�*~�˝H^�YG�L��*w�W|��[�?Yj���DS�VJ�Td`��O"?�~��|�t�(��@U�p�P}P��J��C]����ZL֠)%ׄ�s���`� �>�b���E~//Hw2�/ݨ,�����$+\ �'%*��ֈ_�rꊚ�����/����=L��'��a����	�ʩh���W��|���kTm�9���J&8]��Ȼӛ��	���oX�6c�n��y��1��9��u���΅������V��T�4eW���9zU���ޥ�h������ȳlҴD�Uk;vՑ�ef��	�r��pB"��=��ŵq
A����
.qT�.��^L�9I-Em:��AI$�oxƿ��ҹ����c��D:��;`m '����*��L!r7G�a �ҊA}"��(z?A[��O,�'s��|�b�C��$W�0.	��J����A��l�kk��c=��OJy7s�����$��ߊ��go�S0(-�P�.��Ӳ't�Cچ�H�4I~��`�#ъ�M�XtH/vsE��z筟	����4ߊa߯2R����;3O�����l:>�C�Sc4c�����͕�����۸+ϱ�+�,j	�)S�0c���_1M���I�֭&��|n�XF��+y��ze
xI����;{���Z�t~�ku/�����k v�{���c�:��j�~�HO�ٽ��UO����#8��F>������U���5�q����ƪI)\�Cn�g�z��<�(Ҥ��+6�V���7I;Z����uI&}
���h����g��ӡYr�y�7�8�୉鱇�NBHv6m+�.�J=M�	U`��G&�ͨ^Y�D��M=;���Q�p�d1o�Z�]�c	�W3�3^c�pE�v�J���8��}���i-�]���[�x�B�-�˷��W�T�UX_�밗{���K����Hf�Id]ܶtH!�����V:S�:U�N��������*1��P�!qM��Ϭ� MG�6��Z��MV-#�#%gr���6��[oEQ��*�\����Ra��X��L:HǖȚ�����%nM�u�T�($��D�P{�=�_�[�����}�<[iwh��Lwfn0�0�3�ˉ��ЧN�����* ��\�-/�v(��B�}�8a��F���txQ̝V\�z��gt�Ʈ����H���E4��Si4Ì�\��=�D�������������:i����}�Lq*��j��%o�Ť�Y�ᶚ*0�����O�Ǿ֗� ��۷����쵹����DC�H�ԌF�t+�f|��'�0E�V����;��%��cb&遣��/�m��ȱ���(zwx�S���u���6����(J�:g�Ǻ���7D�G�,�&���mf_�B�ʯ'1�Q����/gI���!t��FtCf��bz��&�+,���aZy ���ÔP�8�����;`A�2��w�ݖI��^�{s�<5 4�Ƚt��&�,���XoQ��q��8�u����f�yZ36`K���ѽ����,�<�A$���h@�S�� @f� ��>���R/����^<�۰�b�?�gқ���GiN�:^��O�����GK7ƫh�`Q54�A/g6v��6Ξ�Wu��g�~��d�%�q��W���i�1��~��Uȵh}�D�π|H_���f\���L�FIN1H/��fU͒#���=���?�^s�5\����qF������j֘��9l0v����bF}%�\�L��'{��y5�-e��\�v�BD^%����S����rDt��(�?�O]�\%4���w��yȧ�IT�㳙zψc�W	�P���D�