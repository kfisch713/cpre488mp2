XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n�Af�'Qm(j�!4��}��R�Q�5=�%�W@��~�&�R\�m5C&��f��hv�k������R��)Y# �f�i��,S��v��4
�I�C<����_Bg�6���y_9�C�.�x�0�e��y�FQ2�Zh%@w��[H�ɹ�_���l,��ݶ ݘ�_�+�rشx�@�'?��W��F{��_cp�|)���u��.���P�tu�YP��$Pa>Jx���L�M���Q�5u����qէzTlK�,�¹�8���H�t�ێƎ��IZ�M������Ґ��y� ��/�����K�{�k5��I�:����K����ȡ���z0���w�a�qZ�\��J;���`�a@
+��:�չZ�S=�%���J�Йm�$4Z��;	=��'O�*�T��D�f�c*�k1P��Ǵj/��3<�e8[#Y���R�%kC-
d���Cb��:����DF����a�W���olH�U7����sc~*��A���z5��A��Ȍ�2ےS�$���Ԫ�TS#G!��������h����;�k<�;}�3mt����^u�1�G���(�2Blj�6�,?繻��������|:���]�S�X�`He�m�N	TaPWՊB�Gˑӆ����^�!�r*�q25�O(�5�cJ����<u�	d��[*��ET]0g!�Y�Y�m��Q- �%�d�Kz��M���Wl�٧3Ҟ�E�>��/HH{�p�hΪc�#(-���f�XlxVHYEB     f9d     6c0�"7�_�Q�euKX���L8���LP�r�O�l�Pǀ�bi�rj�:��[�qZ�E�,�->"b�k���vl]%��3$61,Z~���)ts��:���j��O��Y����%6�~jv�X>\�鶢8n������;��ݡ����c@�tj�e.�g/���c�I�v�3��?�$8��:ʳ�'��Tpd�=i���VM�z�Mb�������\��My���jE5��y�F�W��)�L�_��J����=T��F�y��ə�������Hg���˭������{�NTɆ2��&�Piu���^6����X< �b$˛���^�l�֊�2���|�:m:�>%�A4�)��)��/-�I���a�W��_��͈繦En�6r�aQ�·�+��)K��{� ���o���=|�x�,�n�%8i����s�8r⎮���F�@C|��f@��7��[�Ig `��V�����P�doͧ�t�O�ו�wO\�v��h'��k�9/	��Vpg" ��>�6nC�=&{+J(��*�M+��'� ��8.�
yd�FK�煷�J��"R�$�rwq�	�.u�����%��ϝ�nd��R���s����L�����a�.�X_g�`h����6h�|*��&����t����B���r�Y��Wj�����G�Gֈz,0�Sl?�DF%Iy|_��@��S�;��|�<���H۹9����*��R�����ОO�@l�{�PL�,MEX�r�\}6.c�Ɔ�f>�ۡ�p�u`V� .��n)����O���aV��6��Mk`�Ft���!1��v��9��9��������,����6��Q������N5��?�A�Y�1q!I�f�Z@��H0�,�V^�j�_��P�8�Ѽ��H��B�4ɞ_�`�W�ɜW������~~��y/N|��0A�Lf:�	���*~Yūn�@ 
�������:a.psm�p��Ѝ����/
��u�4�퟾���W`���Y'?]� 5�f�͠J�M(��.]Dlk��ꛈ��W�����D5Rc}|aƁF�Jy ��`厽A?��<���2VA�y����w����v}e�X�����.�#�p��G4����f��T~�b5�E�����������5�E݃��Hu�c�n�@U�� �dj���a���x�0�LB��@@��%qd-z�hIkM51�J�IW�K�z�`��-e]����h0�&��!����� ���
�7f���|�
6oB����� �M��z���>E~_]S+D��i0�+b�BO+S'Rw�[O��-�$@m3�"��`zD��fG�`�G=FR|C����S�TuF�3��t�`^�cf[VKP&�L�n>��C(�i���fA��b-�AO9�CW��
�'%���Qw�����Mُ�6�3"U��d�C��奿�G��b+zw��ɺ^����+�l��]�/�iuu��eu�����}�����}Pv�ć��f}�?�K�D��d�~��胴4ݷ�2��5<�_����U5"ICijauQ5󙌋(�"�&��Z�a
���$�S��)�1i�&���Sc"M�#H�}:��H��Z��������_7A��GGn�;��x�fⓝ2�	fo+XV��қ�1����z&�$Tn\��=�f�{L��΅� d:)����,&v�W��F�!�ΞE��S��