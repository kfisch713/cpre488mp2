XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{�e�-��Vt�X��ՈR����F�*k� ��sL�a5�D�����y�+r�/
�z��a'!���Z-��?�Q���YNȹj�����g���i��wmضg�تZV~��'�ݸS��_��MQ�dB71;b��=%O�9 <k��x���(�������0�~�%����U���_f�������*�Eá���)�٤�Н(s����.�1%�g����t�K��R���s��.բ㴣s�V9%pۓ��=FroЉ��>�ZD�X������+8�Ņ58���-&���l�߃	Ko�8 �N��J��b�pU!���퀻B;,�̏����⬡/Hy��XF	�
kO`]����Elo< 6��><�n���d3ˀ�� ��4
f��i�Ǻ}�9ʬP��s"_��o��8օ��õ&�%�����Ai�3����$�uU��[R��@z�(hF>~퐄��Rx']�&��:^��Ѯ >��ۊ�|�t�/����ɩ�NkF���JӍ�޽^�-<��-�q#��dQ$�.�j�S��y��2M���@7%�/s�˅I/ۓ!���;1f`
����]-r���Iw|��8XX��i% S=2��K�p����(�������j�s��o4Ru���h.��2���k��g�M߉�"T�<>��i�C B��ƍ�o��2Y�3b`�_S�Ֆ����y|�Rh8�z�8S���P�M�5t$� ����.��ԕ��b��'��?��`S�|y����E�u,&zi��s,XlxVHYEB    82c3    1970a��z
�l�p#���J�Ћ<�ԝ6����3�⌏d�N��C���!��9��JN@���O�>�5��ћ�8�wX��b��$7�T��09B���:VI\�y�>Y��\og��._W�.Ei��wx�q���&˾+֋��Z�p���mwD
�SᤢO�~c1�����a1ާLX6l��w(�Z'*adR�&5y햪���ɿt�iF	c
��#�{���.P�Sc�	���A*vz��-u�C2͆D-ahR�Q�p��9�PBI��ѽo���=���^V�E�i��
��B\/U�6���s�Õ`@��<�W!|��&��̦��A���ek�\�=�3qgSNpϲriKAvz�C�^�. !�Q����g��t~��i�[�%ʍ8�����f�;�%~������̰���w�}i|4䎉�o��~b��_Ǒ+�?�_ۋG5]��鐙����U	BI|��������q�5x�)���HE�^8R�y�kp�h$M��E�O7�qRH���l��ߩ���І��D����Fi���~]z�e��i�}cъ3ҿ��o��4,N�@��ro'��²��\uYC{�4��W�R~{��v*�|d{�Ά�Ow��"c}M>���s&���
�-�8�]��1���8�I7L���,�� �l�����g���j}�ó})��+U��L۹��*�rn��{��1��.��}l���fg��s�8�
~�`�{TǠ� 3�HC�m@��k�e��f�or�A��A56�i�h��
��1�S3��,�������uK�`h�I�Q���,E(5߻+�+������'*���f��|@;ን�G���P��[�k�E��W��4O�O
t��XFT��?G_��Ԉ1�n�&Av4sqE������� ΢i��u�]�;�N��2̺[/a�dy6�C{���}�I\�U�q�I��d��,S4�C'�0���wm�ᩜh�� &���*��g2�jۣ�g�(f�.:��	�b�����6.�k��T�N�.Ź%avF�'�c4A�赘����K4��Pb�Kk��>��<����X֌;)7	�,*KJ�1)KƖ4�N\� �=�E~�~���u��Q~>��QqN33�#�oՊNֽ��T�{���f�J;��	39^�%���c��J`���9���9]�����@ӄ셢juv܏X�R���fGL�q��̩�� "ǿ�ړ��6UuO����īV��'-3�|�> ���BT;/��}�������.��י 5ܯ�Z�}�5	8���,_��Ҁ@#*{��-�Zii�C/�T�w �X$�kEX�?F�g}��#ׂ�86�20������w�uba8<z�Ģ:.�X}����u>� �wX3���FK�����ha/��ltW��L�V�ć��$
:L��B5��a�L�s���ִh��l����.Eq��a��h�!�ϣ�o+�@+�� �E��N����?#�"v/,�tOl�+t�.�A]�B��Hԩc4��E�Jb
{�^Jmavi\Qe��alr�2�!$�������'ql`�`����k F�F~vGekH����su�g6|!������z�� �И#�&|��}r�^	�����	��(C��>m��Q��Sh�X�v����V�0G�g�D����$�w�q-�|^�j]�
�^��嚔��2�8�a��@+:Zk�f��\#�
������������Mk��G\kS��e�p�Ԕw���u����U;BX̂#{QD�fV$���{�ҡ�(6��q�����s���z8�"kbf��D��n�t9?�詟{/<��PU!���<�� �&BDr��@�`*�m��{<��b&�}���CSf�.��c�*?�dߣ��^]��Q_��C{0��}���bIo{�Y[��02��!W!�5q�^[v%]�A���f�D0�0r	E@fto�gr�߯EQBb�$�7�61܇��>\�?7����P&��%���_(�z��o&A��"ӂ�f�H�atY���EѮO�-,9�խTd~O�0X>?�_���[����JBsC�����iu�|b\k=��g�3
j_A,�\���C�mZ�p��c�X�
m�%��<&3��N9�b�4��g��}kl��aD^nf��|�idҎ8$o�[���^�9l��ߠѼ=ͥ@������=��ϥr�ɍb_��j�������)�'�������x�ɹ�p͇0�7.фvYD�
����G�c^��X�#�R��Dŕ�ACV�wBej��	���^�̇L���D�1�p	��CMއ��F�8�\�r���RvB��y�m���T���2U�U�/��2�5hx��s�:��J�H�����&���<��V�b	?�Y2�2��������D٘�ȧ��������$���.}<��x��[�	�,.���ߞ�^	�Y�{��f��#�g��m&c��g� ��g����ׅ�-���["Oa,u��#ns�Kޠ�a��WQ���K�Uh�D�1�5�
	����8ۓ��	
�y���3�5��i*@��-�O�����C�Ϧ���,��?�SW�
��i�J@f��1����nI�����/l�;U���I�v���<OQ��w�'4�K�ї� V�����%�(&@�L'�9���(c�Y'�9	ڣ^g��6�1�?Uw�wc�D<Ȯ��Y�`#xS��r�<�Wk�� ����-p��!b�kr�r�L'����6�v�;R����Twv�E���{5�kt�x��$��"	�uj�B�z���±^P�.�~����.~��}J�u�9[�3Y���zT�OǞr����>���(��*�:rf!c���r%�7����Tׁ@)�@�f��8W�2+��p`�4���ScbbA��%p�}����?�����G���R���	X�bZ�撰ϭ+ �i��K�9��衸@�"���׫��R��e��� ��~^��:DD�]W�oƵ�;ρv���
Ŝ�v��.��.>�<���� E&4X���ii�nK�T���'����q*ﺃ:e�_l�e�-̻���X���	��P���J���"g��}��&]hQ����*<tԏ��!l.3�,9u}f:I�8�꺍�1��=V](+-�)H��-��9�_����x����֐O�� v]-�K���v���嘺�J� �t��E��?ћbp�:'����E��B	�����X�+�ۛjXna��߿�W�v|�Ef�����L�|V��BD�H(����B?V�_��቗�u��՟}4��Dml4���tx���
ACA�]�	�0����m{�h|$��uI�g�2k�8b�4u�n\��Ҩ�Bz�Y+�P:M��6��������Vy�L��D��؈�2�G�T�TE�Nyc#r���x�>��e����Ժ���?�C����P�A�T*�FB�,���_��[>���\��t���j�����A4�b��bm�p��U6칣�?D�=��]�ٲG�c���yByv1,ʀ��WI� �$��1.�C.����ALp=�`�+H���\���S���qC��f.{��#�yS�I���=�β�^�x�ɮ��o;���� _ȥ�*�=q(�{��^��	�څA�իr{���y�G��R#��"\�v�Qn�@\H�ɤl{[9Z�
f�=^� �=��j��� w�/�Ti�[��H"5Z����󏲖h��g-��{v%Rs��䀩�"�{/�b-�,�f���WՒ����@����qO��mL�2p�v����,Pi�W��8�Ɋ�p��hgݒ��k���2����ˇ�¯pD�r����&���)�P��ߛĐ���w���~i#�WY��o2�xc�h	����v���I��
h�h�L|�P��ZT�� )5�Ra��=�*�7f��?튺$�P�����Ʒ!�o�>Y�"g��z���`�F�U� ��tu˒�v|�=�*Vp[���xk�M{����k;��.9V�@R3-\s{{�ʁ�a�������8�'�G����f�k����Q��Lk�euT�:�r�^vy�uX�'Wŏ�˃�|�Wp�\'I�/18��� �`�[���r�ޖ9��AzX�W���Twj����/�di��r�!�x�e�C�8^uz=��!��؝R������*b�2��_�b�}�[s�\�=X#�h��L�"�tY�̂�ːu��*$-q����p��	�q��QeT����N��H��-�,)�v�r�B݊@xS�y�?�;����S��e�2hT_c��a9�h�.�1E'���7��_g̍N5���Қ�vC�H�Fɔ��� ���s`{�ڑ?��LSp�aB �y�8Z��DA{#��Do�;��yk��I��K;�>�JD{�/�3L۹EK��f�/f��	�H�  b
0,���,�_�"2����S���A"���i�k�U0��q��)K(�췝��Q��2��� w�/
!�� jϯk��Tx�� [�Q-v�z�߿��SD�֔'�v�S�Y?�yR�Z�Nn]�"�	�
��鴚�U�@!3�U ��wW�'�dτ벗���;�δ��.*�&?�������t���Jl�Ȫ�3�V��5�����W7���VVSi�A����f��}����TJ�E"�W��ޝ@����N�s������Zr�z��f[Q��Lɘh-ӍИk�o.��$��ߔ�Tq�T���G�b�_����Q�u�*�3����ٖ{T�Q�`,(l�P�dO�2>�o8[�Y���D��eL����.f����������<X{v��+y>t�-�<h���F�����)�	��̯B`Ś�Q�����(������'�I{�)0���$|ҫ'����,͔�Q���h��������s{[k�MaǙ�K$�jzo�εg'��?��j�������������$�df�l�͐���B6��8kDSD��^T��Ԧ	�ř��v^�6�_��S��V�5h��� 
 ?��T�+\�����G~1�ʹzD���R4�	;��n�.CF���8]�����b�E���y�vYT�G��Q���>9��Zc��I�����XsN��H\�Ո�N}�� �F븦�tV�|��m�C0Y��K@�r�W�|ZI���g��Q����׀��[���n��49�ʕ	_���"��V˨��t�ac�'ǱI�|�o.����7���.�5�jp)��%wO�~
�l=;�;��ȕ���|4+xg����>�E8�^t�I[P��]�l;u��(Bޜ�������pV
��|O`}%;�*� _	�K�C�f�ܤ6���"�"��n���<oV�篇D^�lj�Ә^�m ���>j^�-��(�J]|e��d�CV���&г�[�H�ǁ�IXNpMA�(­�@Xt95���� )'����1�9}pm�2b,�%�~��0؛�wJ�0g -�^v�98:sU'ѫ}j�B��v	aq��խ22/�� �l#������Yj�-��W"V`%���5�)=�h���2���=�q��Ch�&s1-C9��2� ��5��"����d�83e�����U�h��r*��r� 32��Wb>9��j9!+���MI�5{����� �����n��響��,�z�A�XyAc#h0vjܯ�,���_�ܻzUk9�oX�:���5�-�}����{�f�G����&62�T��J��>���Abźr�ui-MZ�<�cj6REkG����V�����iu�o��ș��L�!Jȓ����Y�7G��q��qڦ��C'j�K� �����2~��"��	^�߿����L����jWȓ�1$�y;u�+�,�'_�j������Q"j����Lf~9����$3�����U��g6V��&Ra�#���)a�d���kY���W	�U�Ԁ��`L�^��x������� �4%ᆛ~��6lqvtz��{�v�G�G�CD����>�2G�����}��{�P�Q`~,��I�i�H9�b�����=����`�P�#��]�>i�x;p��0���걍�T��&FȮ"YCX��ǫ���R�BY;F*֎Զ
��Z!nY��s���MH�P�$,r���Q�t��E7�����j���f��������G
ǡ��ɦ����Ws�4���_�TWk��C`�ud�E� xE�t���e;�'b�߂�fwR	�Q�~�s��O^}b�]�ZØ���w����#bۢj6!jkb���a���N�z�<Zx�pj�����'�W̧O��}e�Dϝ]�Z@��̖N�����!�3g)Ki[���D�HGk�x)����X�{�7��O�L���6ז����Z����#��Ǫ\L