XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m�_�y��0g-��ds�xnQ��0P�:�|.M���7�ŏ'y�X8��a6vo�Q3��|^����lϮr _��%���Ǘ[[�`�M�տ	yj.�,����Ɠ��R3"|�t)���hdw��R�h�ʟs�H+�aȕ^���̑�A �����4��I�٫��s����a�	������R� ����l�ݔׁr�E��y��va$��6h�Hv&�(�O���F$���}Yaf[ݗ�Ds1t�7$&�=����d5˔}�a�����p7�鏇���-9C{�o��D�ETTm.�`��~��yψh�&w�'�[3��O���||O��Qu��	�U`�����b7ƞ�/���qrN`��^u*ܮ��ti��T�v~�/{�jǅ�iH:� �LS&|=S*�}�c5R�����R6|�~��6����b�O>�;��,��7̢|.������]����VTC#ߴ	�������K=)��4�
�1�4�o�|ճE��Є5�(o3��l��p��eU���1?��t:�aM�Ce�F�m�S���25p8�N�QSFu�+�%JA͖0R���@ u�S&�R,u�Ѿ<^�*��h��" CY�R�U:�+m���G�m������c�H~b��܏���E���ay*|[5�c�}D�;u��E]�={�:xi�Q�G���c�;�0#4g�X�d����)݄�,���D[�?�[� ]�=_49(EJ��s�ɰ<3�[X�:(XlxVHYEB    3fdc    11606n�������CH��x]W�L�Й���aU0����% [i�<D�5.�ԟ�*��d#o�C�;)�}:��O�~DF5�"���;#�R�H��(�#�A�ڹj�I>��K�Lݩ�L��Ǉz)��V
�ш ���Kc���W���펩�Hʴ�Ֆ@Ƥ`Dš�h�v�A�Ұ���#8��p��}�6
j���Ux��hg,���7u/�. �*K�m*��%
i�D���j�f�f,�ơ�ݡ*
�=��a����
��ɽ.����ד~���i>���0������:�||�JQM��
��W�4V�^���{-�a�+��m��I,'�$࢝�ER�!����$�P����|M��N��͠\�t��k`�H�_I���s�o�ڏL�{�Q�e���Z|��j"$��]�&x"5�i�r�<6��s�D��kA�������g���e�j�O��H�9g�hh��%�� �k�Њ=Ĵ��������-]���,&��������ν-�7���d���:/t�g�W�����m���pN���y������o�	�@ǨKP��X^��ۗ����6�2�C��}"�״��8�'~��Q�r�M���_����7z]�k-P'��(m���/*r�jTNl��b�0�d5�EvB�n9+m��a�_2���+1[m��a~ɩ��+4�zC���S�/�����6þ
bffc\���^�/����\L,�H��.;8b.�aA�t�s]	�ǻ���.x��k#t��9N��B�F��Q��kL��e�'=�|��G�pm�>���]��������u�^j9���P�q���iyw+*��6ؔ[���|C�9�3�~E�芪ttǊ�)�'��$i1�������8s7Yy��ͩ[y+��q.�|T��-m\�UۑLBM��$ �� �;%��*f��e��2@����h邝3���41�y��'{Q��ͼ�_��'ftd����![2�t�!q7��4�o-�}��&b��ަ�k|r�X���ď�aj4�V;�$�@�T |��&>�MC:�<?O�8-��s���RHVh�'R0+1���]X���V��i����R�"�$���M�R�'�*Uu�<SQ�i1��N=��<e,��6�����~N��<bM�� ����P����&C��������K.��2�cRփ���]��3�ʬ#����-0knO�y. ��J�S�&`�_���{3���^NX���Xwm��HxHtM(�=���[�ߓ�R��bL��Q!rܰ�]˫N͞�����4���&�N�����	��B0�>�)	�]���'����C���g���< +��X���ʅDÊʽ�ж����1���e9���{�5�G~�{2�y%�[Yy��a��m�,�%rb����Mv�wm���;��D�#o�W0��yE#/|Z��Q�����_��p��f��K���¨ZH��Y��>�fIg�5��@%]�k<϶��S��T��~M06��z��K�3JC&w�g�B��?,`����f'(�!޲&���n�V�����$ӈ�Z�vvj��+տ���8Y
5��,=9�����Ƃ���7p������Tx� ����r䷷}�?<��|��ʪ���X!l�����(��� G�k��+	�>���y�j���}��9
(9m�|׆���W��\�������9�!�9�B��:b!��4~�91"E���F�Q�e�OL�7T-�*!DfT�!dW*è8$���\UR�`�Ĕ��A�O2��8�:Gtn��8�\��>��ضHO�u�߲�Pݲ9�3��sK�-,���`�9��/r|���D]����q��������q(3�_@�����*6,��5����6d�qc�bz�'$���a�,�??�
��+V�F�Mf��3���?�L����-���o���-I�0A􊔖p�k�?�ŠNw��n�̲����&����aE��.��E�\�C3��
�?�[Y��O*cO��1�?��m��#�R�g��0��"Pr�.�v��{����q/f�|�� J�t�(~0)i���G ;��>ctv�_[�u#'韝f��A[�G��Æ28a8bN�-�F�e�����}.Q=�^P����C��ɝ<�:%c�D��d���j@W@|���6M��?l�τEhZ m��u��j�px�~��$���}'.�B���~�p���JW�:{ɱ�0�li�&$.�Z��/�v2s���ڲ���$�L( `/Q�7E?*SA7l:��xAF��5Pwl@����kU�f�ōe����˧�R~�	�6f{ʪ��W�G���tS��9�9����x�!���ɢ�+������ {:���?�v���;���� �K�}A%�KV�N%�%��h��m�ԇ��5�w�Y��C�2֜1k'�C�۰�/ڷ��}ɚ���r����Ñ�rbw~1�9LeL���SZ�X�"�~� C�~9.�9�s?���*�N����"�����q J� �+U#�Y�T�W�n;CC�/���:�08sK����Uκ�&����o�p��G�f�%����_�v���؅���`��~.��U�_U�0���E⫓t�ݹ$T4�*E&�!��)�E���w�:]�u������M���J���}���	��}�������-N��r<m
���ťB}�!��6�� ��X.ڻ�{�h<�SG���GM;�pO�ヒ�{�}�No��0�Y�(����lq����Tx��� ��hJ�?=K��
pҰ��sX����B����(��3Âq����{���RN��-���0��:�;��N=C�j̯���{jd�/v�ܝ��'ʡ[v�؅.ᱼd@Ӕ6���ٯ�6v�;d���)�i�j�w퇣�/㲰C��7&��/'�(�S|�'k^`��@b��D�	�'f(" �Z�WH.2��
�ճ�ﶎ$D�S�*�����x����"8��3Љ���0q_l��_���ץ#E}	p�W��4=�Z�5��c����Y�,0��ֹ�L3��K �1�[X�;�!<k��~�7�U'	� &�t�������9ms.�p��\_�Q�_�"�{	��K��s�y�L0�\��6V�q�ɥ��*����#V�uV�m�>6��g@C1�WZ���bjLѹFّ��:f�̡aV�����M�}g�`��huX_�7�eV !%T�&���؄J�Nä�����[K�l�P��"� �F�<yE��	�2"�V9�v��㳚8�����W�8�|�s�Ù�3�N/([*z��pKQr�|���'�?Ihh�R���ߕD�{<0�H��3�cp�M^8�82���LX��O����U+�xO����ܟ���!�sC
0�W�I���z�)����eZ*H���M�Dt� 8��-����}������гx���O�NLvb�����͍kk�՚g=���9�J��4�����R�`+��Z9�c����0^փ���}V��0�=6u�S�Ȋo/E�Z�I��u!�",����j�� Q�
w}����|��B�g5�|�]�o�?<�܁\���k{�{�Ӷ\�m�Ss��{�Um'��w�M�(�V�莗�"�=\����1. 5�+��g�N�!��*�ug	�C}5|)�o����LÂF �}�8 �1^�n)'���W����B�n���������Gt�zߌ�uL���ҙ�@������O]~����O���B�`�F����n)�9���q��|`�=����j5�sG���~��9&�An9ﺿAФ9d Xx�S���vɔ�qG�Q/#�/؜(� s)N& �_�Uf��l����zt�"p��*IJ�TF�G�)�X�0�w���o�H�5jeټw7�򠗐Q��U�~�-�6���9U+*o���r�1�z�!��5�� ��G���8]F6A�Ji^�1_����Tц�T�E�i����j�%fb���ZƱ�{��G�1��=Z���@�H^�`ѿ�j-��uݶ��0����Ĵuf���Llհ掫�e\c�s茀�{�;�6��>��h�ԉ�pe�$HK���T#��R|-�a+�t�]��OZv 2��H�ð��+T_��+$ ����Óȗ�&aԚ{og��|jn���jd���м�r�_�o�oSI�ܣ%k�8��'�����/g1�g��RK�a�fg�s�2W�.�Y���	�өlڵݳ?'v�;ۓ,-�������M$r�m�E	�#x���o�e��[�[��=�}����'���f��Y��2���Uĩ?<]�@�/�yjoʗ�}V`�~'�p��Y	C�ӭ��c{
!��:�0P�y������|�;���_�*!�#�