XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0��!TJ��>�S���{�!��Ȃ1.����*���(�������C;�c"�0�=�Po
����.c��&�3�Ju��F;�2oh���<}�]}����X�l��L��TC�����v+H�XI:�ț+}]L�&�\'	������W+E�`�4k_gv���j6��LY��1��W�.L6�a�Y��cy|A�q���u��1��U�\���4dҗ�Ơ�S;-�	�ŵ�B��r��ֹ_RZ�����&L5VH��ڦi.� yQ�G�D�%x�����j��I�C�=�i�t��r���������u��"m\
?C��kW�T��ngE׍f�ˇ��TZK��~�mT�1��y��h�D�eD��Z��A��h�r��1�Ѐ�f|��O��K�+P������z����3D:�p[�����b�`�6cn��v��u4&?���F\��o5�>郣�vc�dB<I��ف�\��2��v��]����C�4���%Oh�ZB�>�̯��k^j�v.�l�c�4`�жs�ơ�}ೊO����vc(�\��e��x��Ł��d<��tWI��?�0 �e�+$Q5^�8���'z����L|�Ғ�7�Yۦ6�,� т�Y�,�Uw�8�fU������G��7D�[���������b��{U��3�L���r�`Y����^�`X�k��%��#dxxי1��e�BΞg
ݙ���@���4T��1�4n� 1�Z<����
7�;��,�MrXlxVHYEB    6315    1790j����J�������y]�SOc"M�;���5�}��~0wQ̎�7Ȳ���{��yn�O6�%À�	�F��X��oa�.ix�JxZ�C��u3�Cb"��$��9���q�%��o�B{:t/L�n�(�)�~�A���)����'�������s��?��c��23�v>�Z�� pJ��K(߫Y0�r��Ң��@5�xS�H;�	��Q1��#e����,�n�O�����
l/[�~6G$i�hA_�ڋ+K��F���c�j���T}n��<��c�q_~Z��5/]i�u�x���Q3�3hT�c�6E�m+�&}tPN��s	��%@;t��G�A-}�s�|[ʈ�
�˴�0C���z�I�Nv�$����[.ds$R'>����ULQ�\T�X�ʭ5I%�?H�W;�P����͢�?�9��_���g
���
o�z���\]Q�_��� �aa����#nwlؕ��2Z��&Jp�h�e��i�b�A}�j��fcPV���؃��2j@q�K��$[^��#�U��T�ψ@�[	ć�ȁ*_�ROͫXR$�^=o�c��Y��-��c��I~�Q��*�G�l���X��Y�e	�"�=i��[�Ͻ̋��8�l��X4M�N@j�B�׺lҎ1p����K�\c��;��XS��/�%�Vk)�	��Ł=��gK������#�U��g�L1�B΀ah-@�P�պQ>!7'A��	"��	p��.rw�5��v�g�g��(��6����̕���
N�R8/�Ҹ�����`��������M+�� ������`���=���	�8�{���R�<�n���>d��(+-�S���G�G�y��0�qj�G�X0u��b�j&�'~�6M˃�,X1�� ƹ���C�Ҳ���Zv?#��JxCpۢ��1���M�Z�S����0	�h�x@�@a�oi�|��B$c�.�ZH�w|r^���.�Fq!7��?1����P5[�@���+��rFh���@%��(W�HXF�q֌� <��aM�����if�������:T���j�\u>T\�H�f����r+LX�G(C����4n���7&aO(?����h~��k���K�i�s�1��^n)XY(��{9���߻���2����gM�P�lV�o���|��(�뉩�s?����~�����
QZ�\`M���&ڇ�޺�2����l��dK\J�!X-��7�JJz
���4�	h�)ȸ笍�h���������>'=!�̳���cv�S������]:���@��F�2�w�)�X�3^���ܫ,0\/ �H^���e'�y�z��=O��r�_����QU_��Jnp۽��H���S�]H?(t�@o�<��\�DϦo�J�?�i]鸩(��
:G�g�����u2���n\���[�'ʺ.�K}Jt�uy�K!��w�DuVqzY�3�x�Kg��>�4�-[�F'$�`���9�U�	���P�\�����x�,��n8����6r;���3��+�!-�rh%�t�̒�nF���6*R�����\.(�F�%Q����(ں���}�i���-	��?J-|3~���U 5}|Q?'έ�su%��1c	���T>KA_�]X�hq]Ɛ~�	+���m.VM�:$	��{�u�q�0�T75<J�����E�
^�a�k��8/qf:�����5���
׹&�Y�L&6B��i�0��%�Ч�ُ���v�eME��j4{nMG{n����WB�rE��x8���]"���*h�0����&A��J��6sr��*F6g��=V���#L,�݁�ߑ�|E�wDq����������Fs�[�|Uѷ.}c]�g��h�<`WXq�QGhvI��D���V�D+�fH}hI�q��/0��eR-3$���_�֚�� "�G�⒅�3G[��m��sȾZ�#Ix�G/���k���q��5ۼ^!���,鴣-�_s͍k��˾���,59���>�g��XI2Q���t�W�T>_V4y?Y�0\��[>�/ACY_���ѿ��L�q4����Mو�T7/�E�Ȥ�'�@�]{)��$*/1?)q&�R�-3L`Ó�X�̢_;�cͱ��;��:Jk��&��`W�O�D	��x�p�/}�$��Fj��� {F����h8WRS�}�F�_w��\�n��&!4��l�ZO�Lm���������h�@�L�U�~��F��"ؠᑩ�4߾�h�|���E�Ԑ)�����E˙D��^>(^�6����*�"�xcÂa�� ��@�6N��gN��0���k�:u�}u�85�P�G��2k?���dU)P��)U@ޏ���/��S#� �bH�ݵμV�L0�*�������Ě��k՘5��%�`ٸJ*�ۨ5��D���*v���(�Si�I��ڕ��eyp������d����� ?�!Pz�z�4˥'����A�ц�� �p}��!�M#)|]�5�^9jC�̌0���u�]q����3�Q�+y�n���`b�pI�G���g'��v�,�'���C CРc.K���P;]/ǘ�!��*}_g�O�� .=h<	��NI���R�q��M�_����鳹����R����$��zt���+���|k���I�DT��Pyl�n#������>����5tE���'{�� ����I2��9�"l��B��>,�E�_��Z�~[��)�9��VXS�@gc��p/�T1���x��B�Pƽ�>���$��j��V�����0���Ǵ�Qk�0����A��Y;Ѽ�=��8"��
c�@����Ōr�(P��)B�ڮ2>�����W�e�S�4y���y���g��ϭ
���W퀆�Ռ��C����}�@�@?��2�Z6Ƌ����xA/ͅ���}Z��myZipvP�~�Ψ�
��"P��Qf(�ZI
����N����qo馴�6P�B���ݓ'�A�����㸌`U�IXp**-Y�����;c�Ԫm"�3>i%�����3	�;+�s��H8]���TO�c�m��T[���<ZZϮ�h�xXY'͑c,.
`�%(�p)I�ɘc[����oD�ԛ�4A6�.��o�g��DLh��cР�D�{Q���Lj��A���u�Ѹ`H�R�X<U�ۦ��~nSC�R���CQ-���;PwHg��6eJ��m��^$#ɩcM�c�я":� M�y��ڵ�3m�Yq�:Y���}}tIdZIm`�r���-�>:��l�A1NO��^���5IK�ΘN��q�?z%���WR����������P �0���޴�_�@��;�f`|Rb���9���p'�9�W-g�z�z<�0�LTHc�B�ܸ	?�/DŜ�g��Zf��$��G���&�E��9h�#U��5��B��֙�y��v3���'�k�ary����q�I1x@��%I5��e=��l�z�F(���C�J� 3M��f_0A2|���dW�uctr*[
��ΕV"cC���ճ�F�7ɤ�2��滌R�|iL���5��'�	��9 ���Yk�S���¬��L�����Q�/�?�s����E��;Hl��~�]2DsR�*��
�6zX4�E_�\�J������`s�z�Z;7��W?��:���wR����CX�s�J)�PR �b�)��W���e��`1����4i��2ɒ����Ɯ]vkptn�S�hX�n���@m���ʥ�к .��H�����+�%�@}A�@^��\ڈ`Z���^� f���vEe�.ƿSSך�V��5D�HU�Ԇhaf�;�����,Ԥ�3*�[��`5���/���Ѧ~ߛ�(�5瞴)*-S:Ft�2�~�<��P��� �՝0�u���^��h��@�H+�х�1���Y�8�g8iM�+���4�l�Wi����y�x?!�c�Z���1�H�(��畓�D/q�u�Яz0�# � e��pU��9�R3����i
^��x�@R4���O�sy#�Hl����1ˎ�z�''������1?�ðX���4EĹ�P`��[F8x���G�׆�_�W���l��N�U�MF\�X<B>;��ܢ\��;ʀ������`�<v{Ʌ1P�T�O�O�3���n��c���ɋ�M�.���e������a�75n�\����� �T#���E�{B�F�s���A�Go�$�y��c+�r�֤��������=��a4E ��P������c�C
�K���u����o���,��1X�]Ў�qb�*���([�hsD��o�`&k3�j�:����j�$����sg���!D����F�a�D��i���ۿ�Pk&���;�����OAf�<YD�&E{o� {�9�T���2+,=Y�x�S E�I��W���:�o4{�o���r� )�Ϳ��+5�l�}�% ��\R�</������ic6�K�����S����&MlR�}%��0�Zn1���T��m"O�l�ɠ|g����)�������׵B��n�\���j;`%�9=j�+�{15�VA ��-�^^�X+оF��Q�(��(n�Ɲ��B�Q��̡[��S�ЪڐABZjŢY�L�11���$��~�Jd�ʎ;��9%^�>�fy�X]B���[�K� >���	kΰT��"�ch��u�0����,�f�����0�4߿+�Da����'X(�F��3&�����3�Jہ3��,1�W;�˗W'Yq����l�vU�A�����0����T���ř�1^C��=�s�{�;r��OՎ2���Yi���(�}�5�s���&���h���=�>��CĝȓR�,�;k�KVڠ�!_uY%�4:jCC�)3��իip�U:� Y!"�����t�Z�&�iV��j�Nv��wW$
�E�.�f3ƛ�?^�!&�З�^h>��5l@#��M��8����+a�/KŲ���&\Op `;�]�����y��u���(V�R`1�(�=q�WU#n�mAn>]��wv�wK�P�aBj���!=�B-3�SZ���!E�|�±���l�2�<�����%@�^4���!����#:К�C�w�.Ȓ�^�J�Gy���g�u&� �����K�b��㨥}r,PQf��NWw3k���e>��N��E�9�@{�iS�Ivz;i����Rq����K�7C����(�a���U������oPH�dh\�`���Č�v�B�����M�Si�������h6���T����X����@��6������]���z�깳�ۆ���Āo�.�xW��ZaL�NH2�X{;caҎg-�ʉ}�:l�HϬN�Z$m��Z�c`�m���63��qi7$G/�C
h=���o+~���E�z^f
�C�t���p��,�;	%-�0G"'��k��+Q�8�45��-���K+fP�}*2*n��M�z���/�>�WU{T���R)��~H�<�蹜
��ٻI��T6�"茕��=�O���ڊ�U���rяE�Ts?���>.�Y�x����=���-9����o1֏�0r���y��T�J0���i���#H�X�n��3ƞx�4�H7�N��22� =����	��	Y�����:�P�_���Ǳ��x0�#9G��Y��#������O�7�̷h�-n��íȣ����"�M������r=As��UM7v��L���(*�k��=�؜�"- a>�$M�d��u���u0W;3&�D�̢q�^'���Ö��u����:�"���Q��$���2�B7%��_�׬��Yy/�o"Gī?΃<"mL�͎,R̅���	4<1�����P�^a�S���IQ*KN�%� �Ϫ���;%篴#hJ��q�Iq�6��-n���y����*��;�� eD��R�L���g�ݷ�N2�W�D���}�����W��O�`OY8�ˡ-����)�ԣ@,n���ڃ5�R����r�7���9�>��̅����8�h���b�/��B��K���8!`��� a��