XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�]!�.����#��1���O�ܻn�N��g�u3��"�����'�"{��/?�����k��C}xI�o���µ1;j��,� gd���c�0pK�ҳ�
Syv\nޔO���c�Ց}v��M����-�g���,)���� �5lAVH*U�E�#�"�~I*s2ħ����А܆�YY�>녣-�������y�Ⱦ���s0�l�<�1ant������$��[ށ,E�:��bG-�GM?�7�w��`�J�~�@�;UR�̽��S�~�:���ӿ����+m��4ձ��x��
��{��cp�T��"�I�sBX��v���B�Z k#z�z�s�	�{��t��=�îW�5��E��g����'/"�w�H�ڋ��.�[��߆A�=���T�i~���Ì�X�B�E�֌����i�H�m�_S�2u��dGD�b�za��&���e��tr�����Z��R5��T	cL~��9�K<*����15��w��G1ڴ�I�m�5XD�g�X��ߋ���!"w�W��0�x�7�Y�z�6bd՟��sO"F5m�.�|�;\l�yߢ1�nPt��jж�
�y�� T�hkӉ��;`�+��M\aU�%Ý[�X��ݮGpD�7�=H��_�TP��@(X`m)�Z�R�6�W��,l�rҟ�5آC�APT�;4�`��~j܋�μ��y驉�ѽ��I籺�,�Grz�Q?��	�m{(^�PN��;NEKXlxVHYEB    1421     7a0\�?eW|�գd��t�}'+���p�~�l�eQ��<�)�BЬ_o�|f����:+hA�9��p=�*{>t�&2�t��7ڏ��Ȭ�����)mj��gG%���q?pRZW��}��k��m'D���)�8��'��ܪ�l\������ܕ�1�+��m|Ӕ|}~�M���xkAJl��6r��Q)��A�U��)��K�<l�������Ɩ���"�T�mZ���9�yL7�?��y�WGS)b�1Z�<��5��<�Ǳ�6��������o��ೖS�C����XL�1�*c�F�����*���[')ӫS�,!�㦲�5�Q[�cay��!&ʤcW��z��^�5=gx�5�o��5~h�J�3�{����L�2�9d���q#��|E=�<�c��x7sma24m�BE2���"
��Y�|s�3w�L|*�Ϩ%������fnz6��@��xkG�� %=��a�8���9喆�+�f唋��,�bqd,]���|� r�Q����a�
x��Cެ�M�EQ�99�S|�OC����0��J鐼r̧�/q&R��8RɲsB�t���DA8��Iph��'bR���c��)��$���n7E,Q���ر!	/(��%���/�L�d�hv��Gɮ�h��??�Yx�[[�t=�v���.�HP���A��2��ҝ]��iN���3��&f�4�@���y��#z�=P{5��  -ɉ9�nAZ)j�i3U�`�"s�&�����w�vWH����-������	L�P�	�N�(B��x�u��v�<���W܃ �����j� � ֎{���Y�C��v�=ĞӮ6��R����J�$ỿ�̀i%�x���5���;��!˕��{
T���531>裪a#`A�H�C4��tX🥉�1J�4�qc>�@�7���������noX�E+�H7V�����`��V}=8��M����8�,���;�En���	�'�,�uS:L��K1�n�*�`��=��bpUo"��F�aA����m�|��4v&s}0�j��k?�BH�g�t"�7
Q�"׻�~��o�Ш��9�k�i��`b�x�tjd�D�n{�+ʙh
�Ҥ���T��ƕ0������ۭ��~�|-��˸Z)6��z��F�E4��q��=�{��T�SZ)�w��+�j�vӍG��̖��O��;�`H_���S�A!����,٢��-�:Nc��s��,%^`h�$�˺�i��+�q�L�X&��ʊ���(_�"�Zj����`⑹k��ÀW)4�?����7����Xa~X�����V�Ƈ
��?�)����g�rUk<��������n��{��0t���J+^��EU�M�/�F��G�7��~��R��8E/�n~��4Aa�x�=���^����}��U��Q�J��n�c��|�ӓ�@l/R��U���(�x��J��\�9.*���"�v��s3�L�����7tC�I�p�e�/�_�B�I��?gq)���6P�z	��W���b2Y�~:�:� �i�Tbh2���~��U�ںL�R�R��Fs���]�^s�X���B�
w���V�>�ޙoا�MM����;(��5גM��M����a����V��L�M"���CiiU���f���IWu���fS����FL�ƫjE{�����8H�v��m�%��KWDg����HP�gU��BK��������RLt¢�+b�=*vw�i	��0��W��r�_��v���+R�ff�6*��-z��qD�PWV~�O�?b�,t{��<R��8�V��7�|��*4o�xt�'�:U�،�͉�2�����P�
z;�L�����$c���դ���$3:����b|����7G��%��u���j����K9%3|����pd�I5���=�c���