XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����-�3웵�m�CP6�nD��+<n� %0�OS=J�	�[Y���v;��|��ރ��o��`?����!A ��y��V����J8����/Ьk��i��tapڎ=�Y���3>��$��� �)g�_��P�{v��+]�6�}��-�Ʃ��,�@-ܓt�[J�a��K��o�pп�B�U4}�ށ����O;V�%����?�q^�@�9�*��O��͢نO��E#m6�.�Z(j\��V����TV���|��_?f ���,}���`���_���䇗�� cG���8?:T�XX�_[f�-�uL{]����~:�����Akfw�͸N�(�M��\�����2ʾ���Ę�h'a�(�Y'V)��&�Eb�[�La�X��f�E&�nR��Pv�LK�/2�Į��[�Bk|e��kz4������ms�n��4'�q<,>�e�>�2�d��B%x�<S�����xZ�s�ae�� ����q|{���@m�)��3���]���Z�n���ȌEF�b��|x�/��v���'zt��M�#s�m�i�����JcK�M�V-ߵ��_�?�S�y?���^�Rۺ�D���4@-���v"ݲ���t�⥧;Z�u��j�'y��3d$7P�j�0-�6dbT�,d ���I@��q�\[<�b����j�ڎ�Z��3=p��D��_��snZ������f��q�`�ڝ�_�,y��B�%����KfD- �	��XlxVHYEB    3e93    10b0ܾϙ|z��SA��^~A�
��	,"���^��l�z�5G(���t�~��;>3�v����潶+��8b�^̙\��C:�횷��}�N�1�.Iu"�D���P�+:�!�T�t$� �LS¿����I/����^m�w�ؤ��Ed >S�I����.{�Ƈy�����s�$�e�倐H����e�L��E�:u>3ĤD�zCA�l��Q���� ���E�����$ot�j,U]��W��e�X>�X�k�+��a�P�;C�E`�l�C�k8{E��� Z��YbVYZ�� �ZF5ӹ��d/�sJ=����}��زν*�|��ĮԶ.ˀ_ݹڅ�q"�Oٽ�P0��IpX�g�m�O�������3[8+���7�����X#e�ʹ)r��i2{�Y�c�E���"B(66I �sߓ���?n	���Te���*�B5�97��������B ��]'Ytp���K��繞�r�.�� �ݘ����|��#���6�����7Ow9�n��|ʹ�Ӟ�.mC*������� O���'>0˰��л�&�c� �+�}���%y��t�{��jэ�X��i��v?hp��nv����l�f&l�E�tp�֏Z�_\M��FG��i|ߛŃ�'�KI�������	�'"� !c�iX����[ �b9(�N/0Kʜ�a5�+gt��!���~���"yT�}���WVף����c��9���ua�5F���QB����Np�
rqj�l'j*S_�`��R��|5��AZ3�lZ2���uu'Gܩ6����h`Ru,�<Զ'�l���f�����0�9��e��WLQZN�{��R���M��[:��ڴ� ߢ�~%z��;h�3����3cg���K�I�AA��ʭ��>�[7-�T��_�s��w����M˞�=�Jj��N����!��O
��d!��D����k
Y.�:��@��
�^�r��u�;b��ޒH��V�Co�N�wD%��eW�����T�^�E�s���o�_T<��/��Q���-���%�c�G��������r ���Y+{�28W��ϳZ6^�����Q󧤞��*�zP�b%�O�$g���&~�g�r��y[�8�B�E��L��H�K�)n������ �l�*I څ�G{1x�l��~"G���A���#=y��T� �D�y, Á�	����޳*�4_�]nNʢXHu;3�p�� �+����BҺR�����|������p[P`�����Aպc�LTd�=��eã���CS�<𿯔B���η�ا�R��$���2;��r���f��ռ����I�'O��Y>=A������!�C%�,�L��{���hi�"N�o��-ǪDڎ^0uEYҟ43tK<��&G�_lz�X�M*K%�O�$Yn��{���hNW���ӱ�����{���Gےg��=���j�0��V�* L�1-��b;5h���<(��TSao�������|G3�4�3�ͽ����QX�c���IT6�Mo��h�{_3h�=�:��
����!����4� ��X���(k?F�/C09Z�\��!T`]��p��]Y��?�<�nTc���Db�D����a��c=�]���5���1j%�JdXE�J�򁺈�%k����̫�=ʴ��Q@/��3q\��'�b���^�]�b��ƺ'�䧍����׀,�r�:�H��!*�cgeL4ު<#��������u�*O���YC7g8�?@��Ct{��A\���wc�(�������m��%�՜�q�˂��W6XX=v�p�����ȸW�Æ�X4=��gI7fpk��5JaT��Ev��#~������������<{����k���}B�ة���X$�,҆�|��b��$+f)�L�3�3a��R��
^=��M_"-"����)�W&o��eůa�\����#mS�C~i��m��~L�}�?kHCb|iw��md��j��0̱dx|*��m����CH�8c�b�AO:4��y=HU�e�R�/Y�������{�C*~�Fݯ�'�&
u�����|,���<~&2�&�,L9%`������q���$;Cv7#l"e�il������W��`B�_��Y�;Zo'Fሎ^��+��sI==:|y�)�~��P\��X	��o[S&�^�˝S�@�'�a��<]a�H�� ؛��B�Y|ごDNQ���Az$"7+��n�T$�^_�ϤU���5��ሞ����?Z�{��"�	L�!t�{0�\w.u�D�Q�/"�7p]	��ïmvҮOUi&[*�ӯ���Z'��+�k�� ���
[�<��/5�� ���=�憻�\�i�ٖ��!,}Z�pӺ	`9�*T-Y�գ�_W��:`+���ö.|��U��k.jo%#p�s�cR�-9��a��YnC���m���\�6>J�
7��s�b�'ub�f �(�l�7���� �A0}WU�;����e?������`�S��R�F)��@ዄW�p���*��$���OB�oI�8�T��2���*V�ڠ9Ռq�C���2\HzK��o�"�9�{Ii��>>�O����6X+I�������9"�,<���������Tq¤� ���'����� ۄY�T��,�8Tƌjތ�I~�q�D�j�Y�A�~(Xs1��<?��FH�##��)���)��fc����3�{��_e�
|���\�3�|�����K�BZZ%��U�s ����^�Z�2��q��N����Ҕ�} +ں�h?�ac�Y�/C$��1�p�V�F5����O�r��?[z�*'9��W"��{�ڃQ~1i\�]�`�7���k�_B$�l=�2Qn�s�z%$�.�H�m|S�YT7���d��;��8Ț��UUFDn���4�	�c1Oۋ:�N� �*�U�j!̳�fr�s�W�5cb�w�k�����pB�Yv��۬�ö(E�ӯ!��t⨪ߩ(j�={Pe��|(֩MM�"�mG��[J%��u�x��F.�v�R��l~�O�Ӽ�˸s��Ah_ʻ��q1�����j�IW��="�1�Z��>�,D�k��fͬD���0,B69�E����/�T�4�8�t�g���#L��V��b�2����ɶ8���p`<��<2�����)"��졸2L�<�O4HKLݐ\�*½21��Y�䚦bל��I=l'��w��	��t-ʁ�xR=.=D���W����14(�*��?�x>�!9�9���G������Ψ���L��ԔNd�5�l�ȷ��%�X��9� x������ғ#�h(f˸En�#N���ŴHFRьNt`��w�y��|N2� ��'u�1�Δ|���g(�Z(&B��*�������;ے��B�"sAȸ��w�p�Bˤ�xjM|��Z�4��RI��]Z�at�\�u
�E���a�
��Ou����i!���G�2-�C=��x T�c���mo �%�E��l(�y�.	y~�� �PƉUy����\��  %��sX7p8[�{	�� ��z1i���M\p�d��H�|2�p�l��E����o�{T\����k��e��k���҆P�H&��U�к]SP`u����7��9�tF&��}�������̩n���1i%
+t���ϪB��W��+m��{�:
#я��/�����
&.�k� :��}:9�
��4��~����7u-��"�*���ver۳q[6,�����H؝w����2�n�e�kB�Y��贻�W�#n`�a��	���cf�S�9���L����߳�i���!��R���<���H��!��޺	�姺�����t/��O�
�E[��M2!F\����$�ǁ+�#=��:��	��`�slKc��I���<W�Lo�4콑g����Sk��j����>�8�=�ؒ�2�_臸%&B��+��آ��B���9����ʛ��q&�S,�>��|��_λ����/=�'ȧ)O�k���-��w���;��_^�m���+(N�|`����F
�H<��mk�U&=XgZ���~.�	ᴚg�C?�c����t{�S�^9C�pw1,)3���<cOM��K¼���!��y`�ؽ�\�t�t���Grr�^eO]�/QO�G,*��CcG;�Nƭ�����ڊ�