XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������H�<��i�����z�h�?R�c���,�G�s����k�ϑ������?�c�v;��+y�4J��-�R��v�7�Z-Qh���#�DLw7��?3s�}�������$piK;'����=��[�*Ѧ���T�o���0��� �� /�'D���x�b��H6]��˧n��b̽_c�� w(Dn��3e99��~�����"ٮԉP�t��)�{7zx�R)1����_�lC��ϫ0�t��쥑 ڏ�fhs=H�6!�B8�,ɧ`Z\���xM#`d{��.$���X���wl����%�Q#���b��Z<Y�*ye�O}��}A���EQ��S�2\�O�=���R��d[������b8d"��rZ}���W��Ș�y,B!�R�!k̫C+�'���ϻ��u�~s	�Y#Z�h^F��D�N�r,�){q�u����iډ��P�Ȱ�������[�2V�Ȃ�L�2G�}㺠nǘӷV����p�<(ĹH��S�5�km0��h��5�!��Dw�i�#��))��|����~�`���KT�;�s��޳i?E��|���}���2�c�l��TG��J�)/��c;����7�U���k:����Dg�L��n�3[�ܸ��7����L&�Ů�ډ�eOs���ۭ+�#��+v��Ǆ�Oe�B4�Xފ�x��q���B��q�p�.e�G�&k9O�>�c������*4X0�]%����<w��|H�M��^��iRON�An�Q�rFQrXlxVHYEB    1ea4     920��bչ��?�揈4���]���}H�ى:��)b���_kD/M�Yĭ(�y��/�ܐ)���qV�s�ʄ��E�a���d��{�q߷�r�����L�l��~�l�k��dn����QȤkG�����f�3:wԙ?qX�g�b��ⴈ�\(�PJ-�,y��Vت�dЋ%�zo
���WW~��zS9�c� 7 ~y> Ek��$n�{��4��&!�5Ҟ@���O4B��o� 춘��Z8xS,k%�&�bQIcsv��D�U��u�i��-40��B��1�t��e�]矇��9��|9�rF|���7���qM�8� d��5s
���׍�¢n��I�tN\ ��A[�{&+��B4�n5��ݛ@Y*�y�s\��V�2�H�S5
�\F֦5V��~�_{�f�y{��$�HV͡�:}����6X!��`�c��`��~nw�o�M�H�s�?��D����
���~�p�aA��;����]wդ�  z��r~;�)bY�a��[���91=��Ua@`Qa�8�����L���E8) 0�	[/h_� ��z�Z,�U
�L��i����������I,w��~�f�k�5��<�����c�a�8N�ף�=��4�(���0\Nly����8d��Hx��q���T��JA�B�b��{t�2M�ng���99�z����t�؃hFX��#W��In;�/����Z0�՛���r��@�u��~����䡰���[�o���V�P&��|o����|,�!�|é�!��������g��8ŉ�7����%2Җ��Q��`�dW�����LY^Zue�i'�	�!Ћ=�R��W�l��Ӭ����8�sdF���i�l;��	����E:j�]d�}Ұ��x�y���jqe���Y���.X22i��)x
�%s��z���#.��,��x��N���d������<R��9�C���-+m-��m#3�%�޵��~���3��T�Tv^+��n{d+z��,{�(�"��	����F��a<@ߥëv����40R�$��bQw���"bQ��JOc�S�p�g8��D�ڹi�r��'Om ~yRת���'��̓+D !y΢V�pc�Še(�4M�n���gΎ��|8�j����MC=�{�^=��`cT�*��U��z�`�@d	���t��������A��\�*��6u��� �.�y�bK̵�_+䧋QS��J8���K��]�����Aw�(� �6��n���)��屰f8�[��8���������J�B8֚u�I����vZB;����0��C�����gw2�<򿿐�n�Գ���4ޱl���$Xy�\��IWd�a�Xa%L83��Dp�>�r�R�z�%�V�=��+�R:|<�W���Y�� ^Q��f�Y��К��KR��!�����8�T�o	�耂0
�[�7�o@�ڜ��Q���P�tt�f4M�h��@���i&[�$�����P��AR�G�;}�|	By��pUy�a����#�~��c����o�g���5���E����}����@D�\�2�U}�Z��T5Ry+�z1b��IkK�g2���-\�q
k�����5(��g2�/��:�/a2�k'���h��a�I��0�m��#V�˷!���yLL<mQC�=�Q�pS��Rc���Y� Y��\�\�~Ss(۔���c	��Ƨd+��y��Ѥ��so�7�@`J���/F�9��"�z�'��y�yJ=��
h拄�0b��!��E�����-e@�Q�����ؼ6D@��N�@>ɸ6�G{��i^�A��ȠgƐ�w�w�o�Js�0���J�R��	圊ս�I���>zа����\�Vh��.�qKj�[m0N�*�_�	�r�zwJ쿍2\	A/t�V�[�Y`I��
�L�v���{6����c�1���IX([�g�s��;:]�Ta�m�y-��2nb[���nM<D̕P.3|@���
��_�o=H�V���$�ޡR�!��S��ݛE��`C��4:섂�"`c�ۥ��1��w.n2�tW_^�q.q35���T�a�S-6��u
+:|����y1�H9$J���h�B��dE���!�|a��a�A�d,���;���_�!���|E�D�7�i��]Q#���Rfa�"��Ə����}~k��{b�N([�u�PWe�"�F�9(��M�)S���!#q��2fI�@t AA�������f��Pq��4Ws��j��΄Y�Gο¥���K�ھVӃ<x<(�`�d�{]`�������DbO�o	�r#