XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x:+�F4�u� %5tƬ�7!n�� �/��S��UX�WK����v�oCF	��QH�W��NY�6��X��&�qfM�y׀��lv�Rͪ>O?�������o�CJ�C��n/q���E�
Y�E���B�f�}����Sܫ:�8rxS��O�쮹����� 3�/�O�y��E:X`�'���Ix�Yڐ�E�<���Sv�n�w�y
kc��<k�οo��}�X�A@��#�쬤��K�8`�u���{+����nfx)��ЕSegG;v��w�I>���������T���j�����8��bˑu%�=���H��nC��]f�Ӂ$�bf�0IjO� �n�^CPibz@k_��>A��a0F�Sh�z���#�u�Yu�"�����h�S>	L�"ǌfY���vY�]��K؅e,��ħ���O����⣿h�q4u@1��+�$ZY�>��(�����ձ�x���<6�I�p�υ�=�Z�91�G�AW}�(�@���
����L�D��Zq�*����2yl���6s�l>a~�}�i�i ��.Z����b��/��¯6���}�o�`0� �<L��।��2��0��s8{&tBe0�w�An�
g�e�|�M�(�GF2/_t$����'р�^��l\S�@�*�pKY�b��-�O-A��[^}kØ�����qM?��U��OK�d�t�f�ܭ��8:�X?�a+�*�6UXlxVHYEB    4284    1110r���`2C���4��$:{��w+�Dz��k���,�WC�a8�ɷW�Q��"b�)H)��R�_�48�,�/������J���%p�ڠvV�$�ٛ�]3�o��d{R��q�|7�MQ�\N����w�`1(�B�o�H_��9Z�*�_3���ϳ�aޝ���/����bm�C�$�U����Y{�x'�Y�1���mP�p�a��ц�c&[_+�@�>"G�v#����C�5��?/���[ ���������)e�0��M^��%Q���
�k�����	�G���Uz�~Z��hE�yS[��ϭ��4Y��f�g}�Ji�����b���-0�_��A\+���_����"l�@���R�pA��W���^m�1��;�7��F����d �>6Z\F���F$�x�$#�{���Q<��u�F }ʟ�<İ/G+a���r��O���\��e���03�R����,
�@ c�����b���ˆU=��d6-,�D�;�4��&4�'Y�3ґ	�;qI[�:l��3�y���F��i��.;���{���{D�
u������EB�+���q�6��#��[��l��\�#��)�Y�Xs��dVu-�:pT�Č���I��|;"n�������Ulj��3��D������d�U�DZݩ�OO�k��tTΆ�ˆ���]��Ȯq
Ҡψ�VM�ǔ)��!z�A-��۹Jʮb��5Y��hd#�� ���X�a+���£+9��s����Hb��e��_/��w!���j`��a"\��G�ē�"��
z)#躮�U^M�gs2�+[>A���\�|���T.~	��Q���7��,��`<��w�ൊX.?���]���Q��2۽Н<�
�������*D�6Q���7AFP_���`�H�?5��	K��"#�gq4o��ܥ���h&��.��w�@���E��D	?dB�"#zx���SL�*���LA��)i��B�ީ:^��_;���u��o:^Z�������t�����d�A����,���{@
���@�9��?Bm��I�8�E�)lg:��4���5��	�,W�M�p\{L\p�8��PjM�3��)����!��C�,��T�P�A��3V��kܰ͌7���_�GY�{�����9^�nB`|���Cy0��ߗ�f�����4� ���Y�i^�F9"�CM����b��tؐ �h�%�����*N8R�VC� V+M�D�0����q1E�s��;g�<T�[��X��|����?��0�q����v��\G�X���e�rd��Z��&��t����%Q��X�}yr��I�|o�P0j���������3jK�1�yd��x�6|�aF����x��#2�����1lnڤ��b^��j�����`�����O����GT��0���1ra�(�]J��|�zu_������=�W��(�l�|3$��V���P�fŪ�����,��YG�(�0�wX� �jս&x��JbuЫn-*6 ��v4���R���p��^�*��F:D��Em/���\Ix��׈���/�B�M]�E<ո{o���q������Dve�x�O���ѲaF��[�āk�hj>��i(F��ܧ��{��4���C�06�n��Q�+vG�h��H�K���!����m(C��hFT��c7%�EL�T�/֐k`4q��>�?��	l����@jrd����K��
9A5[��,�j�O�5�)<?�Ǹ�h(n�9��mY� �]I)o��I�����p�ve%ܴ����9?��a�Sls�+dGqK�f����ٽF�ρ�����ʙ�kw"���=җ(��6�oz�q��V�,������K.��6��g푩�~��ÞUv[����2b�REFJu[��S�ŎCӋ�A�Q �{B���o���X��h��ik���1q�m��ƙjvi>���tN�+8��V"�ej,���Q��X�v}�t���.�-�-�K}i��tm
�7h�_	�b�@��BA�������HҸ^Ӄg�,��46L 6�^9�=�� ��t�i�-[���|�K���N���	� �c�
tNQ���ĻS��t"� �/-��uc�UNx��	������{A��ΠD�����0���F�������F[-��P�a@~�]��lC��܂��w������-`��Ape���+�'Eb�UB��������cB�*EO��(��W�{'⩒C�a�Xɴ{&�vۍ/9y��_5�n@ M�fG�Ӫw�w(X��O�ȼ�]����޶U ��7VD�!m��>YUcM��{%y��uZi��o����l[n�����ʵf����6Q�#���頵�Ԭګ3w4�8��9��|�Ǿ=P�u�᧰r�H����m�̜N�ϗ�8���(�K�xr>{�%�a�e�P�8Q1�Zt\��O���	��}o�^u'f�ˬ�Vc3�}5�M:��%/PZ�đ�jbX̷*΍Mȉ@����q��תJ�Z���\���Wmw�J29 W����XX�v�I�q�bh�,V��v4��,�&�>�s�@T� )`�W�ِ��A��o�CD+gr.�&RbK�)&����:�����|V� Ă�W�'2�ˈ
��oh�r�ZI씯NmF�g#n��Ťj��AC��)�����/3~8țHo�K��4S���]iT�����5i��ǎ����"W3Cf��_��x��u��@f]G�@�&8A���̣��wM��`ĺ�@K�i�$�XA���3����H����'�M�W�s�6�lL2�G�#:&���`l<4X�H��x�"�R�@�߱���$�n|j�[�H�_���#��Wų1���m\����Z}��7f�:��2�[;�w.S��`dԃ�Ħ"�+Sgz{�%�����v�� pT@�~>�n�k��|�v�mz�=7�?2x�7s��&�(����xV��hp\6���_�d�W�:!��t�RB��"^]̮E^@��i��/߂w���z@2"(U���\Z9�_����+,%��af�E�I����Ԗ����u�_c"�!�M�I7O���� r��©BT��W5��gp���Az۔�>��sI�Z��ZV��3������׳���l�x(,la4�dZjյ��.��w=���1"6�j�T����U����i����6M ���g0T(�/���ZG���,P������v$��9 �\�N�3��?C��`�R���4�8�����,,�]��������|͋������B��t'���e�F�.���s-0C� ���{iZ�(& �ͤ.�2zY��a6��ލ���߹����j����[�^طu��Q��M���ܷ(ħ���㿄�ߩK"HϢ���e`�~w�V����Lw�W��l3��-�)���
�7������������#�Xz��)�Y��(/����i:�}～KP����?mw�����j�6�n2x+�'2y�J�S�j)C���i���'C��9�F|D�`�A/w����Yf��B�ʷ1�fQ�}�������O���
_��6�Q������q���V���b�	�& �;�m�2���2��&���R�N��T�����Jx�[�J�O/�AYOY�o%���6�v����XDO�;������������P+��v�>*F)'.2\��wI2�Cq�J�%ɘ��u�C���-��C�BvM�C�Ԭc|6�wC�9�� F��͔���-QԼ9M����6h�3�R2=�+R���Œ)3[�K��A�'���Qm� JX:xK����ތJG�����;�_N���3Bv�Y�F�W���1_(<J�r6X�[n����B᳥��\�8���Q�PX54�M�T9����Hm�\=����ߐ�;��Nsks6�J$?=���kuCQ�8z�������A݇��'9�ȳ���ѣ��L	/�rՎ��,b9�~�]�ѤzV>�h�TJ�k6�s�L�);�B<>yO� ^G����Ws�o�to��BP5�hyx�%�7�-��~t����5�H���S��F%�"°'��!��.i�L�k��6|rzG�u���#��k��*rOI=��FV,xU}��j�{T����-���7�|�g�0�hb&	�RK��t����=�[gׅ���t%�GK��u9���0m�zN�6�o�<M����2G$�n��ә��:�Ҁ7 �}�+v�0ɆϴFSS��%�U�
�R7���n���3Z�����Bwҧ��M���`����GNfp