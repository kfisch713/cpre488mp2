XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]��w�Ŷ��BLW^�J����@����_��%@�[[xLP&��߀��+ɍ04M gL%»��</���+F���󣢃�F��)!�BF�G��i%��.���򕣘��[����BL�P���O�/k��6��V��(t����G�]%�:绗�&�V��*��/��y�������H� y]V�6�"�뽑U�st���`�f�E5Q�{?���M��`�[~	��B��?�*Uq�nH&C�
cc�׌.��En���3wz`���g�F�],�_d�s㯸N�?������Ǘrj�����f��M"�n���@A�.
�����Or0h���|���g���}:ʈ��Sj��I'[��:��j�i�؍��߲3a�m:�S��� $�C��/i�2��^�d����Hў�����=�]w����
Ϝ�{5_�9�=�f��3��:so ݻG}=|�`g�,R]?Mŋ8=Y�p�')B�����8�L=��<���oɼn�2����� �S�.@6a��E��R�led�u�(r�k���t��L[�*�b�)���.}�>��#��G��@��ŞHeB�̷�z��KZ�}-��^������Z�))^��y�T�9M�\?&�]]��H���G{.H�:\�yӐ��r�^T*m�,~"X��sw,��S������6Vh�����ǝV�8��:��K����Y�I:RR�8ٌ�L��\��7��S�+��Bu�.A��v�b���P�I�WQ�<%�XlxVHYEB    2892     bc0�eh��NWٵ�n��Tz�u�����ydx!_Y�]�a�)~. F�&���[���Q�t&�p�	���'x�MF\TQ\ܙ\ga�@-{�A���t�C&bb
П�0�?��f�@p"���P����[�`t�M��i;���{G[ʡ/^��Siu*_ʿ�b$]���| ��4(��	�����c�}@��-���s��G�7�ya�΋���$e"d9X:(��W���2���<�o�O�)���'#D��<���n��d���Fȿ��>Z)��!�)�[�V칑�R���Qyh������{R*`������-��&C���k�Vr��ɂ��ٛ�r{D'N|�4���6XoD���F2Y������'.���lͅ���yZVO��YUa �<�7���v�����(��	UЈ��%jmY(L�$ӓ�-�~ks��1$������p�W �9�����\;��o�j�q�� �����K�dY}+�Y�.D�4Sٖ֨�L�
0�U�=u�a:Jt��O�CnlD��
j�cл�i�[6F����Po�$�&�d��W"_m��NҴឍ/�H����%��o� Ţ�kG����ZjlѤz?A���e~��k�Ҩ�� ��-]�vk��ѕ	Ai�\K:���2��:��þS�c�(�����jR�ݝ�8��j�'cH4�]����p]�,��]Bzx�cM��Q!�nӚo��/~Xb㫤��]�Z���yN�SE�s�k5 �Y��IXp��0L��Tz�Hl�"<�L�
�8Y���@}������H$��c�Ow�����U^7��]a��k�6�eȧL�A�߷,u�m���c=t����L
ʆ��6�^����Й߁���hǒF֙e(F�� �,*0��m�p�|�[[��bеy �^��z�qQ����gh鞝JC�,�&G�VY@��g[��ߏ~C�t:q�	8��\/8z]N��b����[C�V�y@ی]L�j��lI�@Z��^=��K�SBj�@�s�bzs�NG��uͿE�����F���׃J��ߩx�kݍR�a�[�-��
5WEEhR���$9ұO�C�$^���l!��,E�@tS� ý�(U��)�nJ^c�����G�7�CUΗ9��K��6�g��H'�U��w{��w�1/��{�����w3W����@��)�� L���ㅾg�[��N���à�T�lw�i��ۂ�Y�ʪ����O��o)��y'	�#x��n-�"�F8iB/����<#�N���
�,�_TlԦu��Ҧ���媙U?�ّ72�X��`gy+H�G����0ߍEW��m�px�N/� D����t>i�����Z����G�r��x��M���	��� ���5O�N��L���i^�i�t��H�,,+a�e&x6���j��,��7�2�Ajxu2� 9Gm��¢���l�~ub�Q��'��T��C����Ii����ʼ��k�����FӍ}�M�G4��x`��Y���A�q<l��E�_�W^jw��]{%���W�Hc	�5�CP98��!���c4q�B�"冗L$>����fY��x.�G�/�ʼ��n��
���`��|p�Ƭr�N��l�|8��wC.@33�4��?����'�������?q�x>���"YS��g �Pvx��k�N� �%/�p �B�[C�����:�BT��y�K� �@�SD�Yf��og��%	P��p��ʜ$�U���
<zErVX����ɸ��En�%%q�Te���Y���#��㵔�o�n�-
�RmJ?<�=(�l���Bp��+�#
L��-$A�~щ�*��6�9 �����޺u-���-ɤWu�"���{/-�2���������Bf"F��"�L\�vlX���Du.��K�>)�>���Ȋhdl����Xj��1���;��s���:�'�O��Fk������zn{?{-)��7._��:e�~�z�����9�0N+AMHV�[O����QND�]P�.C��C�HJ�r�q$��DY�-yr��29|��$]/�!�-�%z�|��Z��N�6�e�����a��w�c �IQ�ʒ5tKqS��pmM��iuu�Ɇ�%�J9�X2$��9�9I��zy.kMD�;���jX�!CQ�,t��$�G����F y��f>U '-,�9�W����JoyPμpe��w�8*���^L�9$s���V_'���˻n���6�@xz�&�&fH�`D�A }��$G�"{�#ⷮ��s�w���*X���<=��]$�}���4�g��pwE{/��-�֥�!bI.	�R!j�G��R��3F�\ϲ����4�_���F�7��tp
�b4��A���X���ձ�������~X�M��t� W�V��^��ܭ-<�v���m�NB�ʺ:�{;��L�8��w���!���m��q�JnX|z�ƺ�P)�8��.sG������I�����}D'�-4�u��7�藕R�7�*�<��7j���re��zĕ��e��Ƥ��;!U�λ&uo>��g�pR�$�nmV�C�ZId��?�(�靳gC�4BgJ�2yxQCʉ��^�������*$�����A�K�^r��%�B��m$`��Ir[��8a �;sAz���u����Q�O�����JF���@���,4�;�|!fn��IW�g� ���=�^�e��u�8f����LoR�=I�w@K����5�Y�Kh����B�O
�@ڍe�y��x�	A��f���:�r�8���_�����a_T3��Vd��$�����[-e����	`�T��wRT��������_=\A,�EEʒ����I}'
/{3+����=W�� ϻɔ�ػ����  �S��ߘ�l2����Z%y���ǿؿ�a[,�����`�����tmâ��Xaƴ7//�fM�Pڌ�4Ĭ�6�7��_�k&&;,�h+J�?�	דֵ�