XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|7R�!���@&Qy�T��$��j�c?����C�*9����V�$���QJ���=^?�bKs<�9�hJ���P �s8��Q]�<��!0N�܈j�X�wuW`ĕN�2��%���fj �%���fU�n`�w�U����m[d8��a��]�$�z�
^�O�XI	T��6SC�/�;.n+��yc>�:.?���[��`���~-�L�.�L]:���3D��}�b�����7�j�xoK'���=zѼb�n���-3�̑��"����T"O�o\��X-#"���vP=|�]I� �n6��v��pFd���v�psX4�P�a{�Q-�P�uQjL�*�XſK;v��"�{����D%Oz� �_đc��8�9�2s,�f�G��n����B��QW�)e&؞E�hhOU��&��o57	-�=
�L�-��F�?�@,��������k7ue�� �RK��
��IN��d�QXHA��xF���;�Y�VӁ�b���.�y1�L�޽�e��$��T�y��������bZq��5���F;��
��CQ�ԙ��Wf`^k���9]��h����@!%Bӛ��{ta�����]��F�Խ�6Չ,l�)A���NV�����]O�Js�KM�!d\I#�l��z�����ep�	��e�亣�3��m��_��㚧bd�p֫�8�*���zS?����f�w��t�84����0/:c �}�2�����'8��u��ʸXlxVHYEB    70a6     b90�(�Z`s��Մj�>�Nz�	"7_��B,aQ������.,yj�v���G0��(������	8-rC�e>�Ԕ��*�gZŎ��!����O�8̊]�,�&��x��+��>�<N�.ɮ2H��AR1�nh����UA�JC̫�@�_�=�	6�㸖p\Q�Y��z(�-�����~ޢ/��}[� �ь��4�BE��)��ʉ����I�k�I�TW���b�s뻚��DD�'�+�����aV>5s���7 �f#!,#h��8G�8i��p���
t(�JK2����۫ҁ�Gʹ�+�Q�:�&gń9�!X�Ch���ꦾ��S�mυO2V`�����S׷-��2Mt��1�h�,�fehl�O.�}�*�,O#�-�~մ�زT��\HV���4��X��y�<�g=l&]�[�P��D�ǑŮ��C�O#��w���b�\,-LĀ;J\���>,o�m��� d����(��O��v+#��(O�M�(�CQ ��pqLt9�I��	���4B�>��|�/V�uj�&O� �}]���s�3�!k5� n&�%��Jį��ց6\AN�>��s��Ėwn�#&P�+���y�J�ٝ��Ϩب(��$���e��V9Q�i0�_�{}cC��L�0�1�C�ͻѤ|�$x^���m��GtH7����+�4��qR������cm���"�V��(�d��Ղ��}��-u@Gae���W�53�,H=�0i����6�ˏ{��b|}1�?�ed�{CS���CD��ՄD-}��g��LU\��y�P�B%�E�ԯ��v؇�F����G}j,�,�\�$�I���C�bb�_�ǿ�=����*�=v������G"��5QD~r�A����ӈ���J������z)��X��5C7q��4��"�gopE�x������/2�*���ޏ�G}}2�;٨G�A��>+f���.&�nZ��)�5�f�f�r��Y�r"Q�H� {�K}HH�!�� s�'�GM}��o��,�0ǡV��Tv�)��ΑUGm6Ȳ�&�|*���ZT.Y�N�ѰN��3J���d�לr��{�����|���a&d��!��[`]4���51�����[��g�kJ`� ��M�����@�\֚�a���ǭ0+�s��Vt����.'X�-]v�8rUw�ψ4=.�7�|���G�~&�+�^�=:	�9�O�@�z��D1p6���m:z ;�hQ�ˌYJ�&���8BI���O�	�%^0(A�6sQ4I�r
�XcL�Bv�k�8K� x �J���:C]��?Zi�4��-M9��s�o��8~��=���]�����i�����TQ��S��Ķ*1���&*	4�+#�2�|���N�
`��9��V89#�@�s�ѽʙ/6:�+��E��Z���õc�*�`�)3�C�\�;��JͰ���Q�=^��� wA�Zg�0i����q	3�g�U��͖� �������
�R����/�,�W�Sͱ��j�;T���������dZ��OA�dZ� �x#v}8P�nj�R@��((�Я�����2\���f��ܫ��޸����H_�N˟{�q���w�~8.j�"�5����j�2�v��5�._cwm��s�Ώ Z�pu޾'��ߝlY��c]V�G�f��mU_�{�\��ަ�`����������X�G'��A��Y��$�H=ʆ\l�Z��H�p�-� �p�$朝|��|�.����3��C�{i:�)	��r��y���2����~Jv��Y�R\v,K ǃ�h_����������,y����"���y�#D��3���`|�y�H��B�RYR�^@�'֑�:	�����d�n�9U�n�l�专Q[A-P"y���]�VdX���K��:H���%�EF�k��[)
�s���i���x�?' 4�~\Á�\�J.O~o%\S�.y ���&�Isv"��<o���b�e��Lj��4�S��es6��"��L�A�-z�9�nK�Q!������sb��MP�`����'��q�ơTH�I�*��֞V�r�����+|ѢT���髆Rg�b�>�ou��c!�����L7jv����ǮU���J�e�h�mn�!.�������z�iiA�nh!�%-���� ��n_���-�I�8�{k������/9GR���B�����0�<���*���X�5��U�S+A�7�5in�ջ��~�=���л�	�@����ė��cMz�q���hJX!;�8�=*���L�`�aĲ��fO�I�d��jk��v�8e\��b��N�W���<y�&��#��5E��AI�7[�((e�Xm�C`�j|��A�e:�.�=B�M��*�V�ҥ6^tn�Q}��V8�y)<�(w�Z�1���0|-�#�
vC�36��f���3,a�MzWzG�����o�fė`�l3ȸ5k ��? �6��"�.�,���; >�$}�78�4�s��A8~!�	�i�w�B)�W��ܰټ�ե�5��<|y<���T�M�!�_�!ջ�kl�<�î�#��	��K�"��Sg�����G��Z*{M=^�\�Y>y�do���oǎ[���_\Gm�ɱ:#r-����˵MDJQ	_�.#*�Rw�M0��憤O��5�["�,��i��f��<�*T�/�^@�	��Xj���S�����{Y�E>���L��y�L�qr�C����i�!���k��)8�����!��"����a�%�gt��r���������h����B|3L�Q��"�1>o=�	V/��g�_�K)��ߞl��%F���\��cƂõ�2K�tG6a�u�q����Y1#!wAoߖ]t@�~v%��A�V#����Tc�E��v�|��,Q�Z�����}S�XG���]b/