XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��m8��U�k��8���sgo��u�U֤��R�%�p�䋁NVts
fL��f`)�����H)��
�M�,�@�B��[��������hkhM �A���mw�\�����5K����[����u�����O��0X��sJC3>1>�㥙��Egfz�����_�lo�%�i�;�ѹ .����1�&�4(G&�I��SX�9p�R�D�2��e䦧�$���@�	6�6R��Q�;��v @Ӵ`K�!�?_�>	�`�bp,������{��et1W�Y�n�
�Z�����>�T�R�n�#@uq{��DB%y��,��zn3��vTqIE^H&xkCɳuY��Ĝ����Ch���-eA�^ɧ�Л�?ɔ�~����;+Z�0�O2%�J��$�1�Z$I���T2�옒F�C����d<ĸԟ����aA�|���Om�r��Y?~�V��t����C4r/��a�i(��Tr�&��J'QI��+J�z������k^w��M��N�a �k��V�}����*!��^3�1S 1Z�\�(ȇ���i�P�-zh�������U��.�eK��?����m�w�N���$'Ҙ�N�5FNK���:'���I
����ʀpR��B^|�D9Rch|��缟J���!�����c���$1�U�[�7`=e�np��v�����|�)�H��@)�fKn�,�{;K��Lz�.3f��G[�u����A%��#H��בc�x�e��f7A<<�XlxVHYEB    3fdc    1160�ݜ�Rv'z�3�n)��k\=$,���ͩ[�4Ԏ�R�� ���N$FFL�I�*`��tn*�!`�_��/5�ui#Ul�`y��������[S-p!Q��b��W$g�@ �ܺ98z��D<��no3�rӏ)�����`+���Ks�GЊ�cF6�"YN\���U�?���"�S�]F����f�Z�,u#uD��p����W�V�_��r��Z�y������÷��f
���(7X���fA��(�n��Ve���oM�R�JɊ��5?����H1�<W~��iT$��7��z�ɳ� |QU�#՘5����,M�q���E����%���?�����3��c}2��8��v�hE����]U�Ÿ\�i��M@t�����f�\L�C�JL/���#�{|񐕻�AC�#!��}�C����y��b�i+�w&��	s0��$�yC�b�Bz٠�u�"�l�}u�x����O�OCfu��4ͭEÔE�`��\�,v}�m��>8q��I'}D\�Rzs�)~Ppz��Gz\Z����6�1��r�H�eȑ��*2Ixh�Q�� �R�6@#�z�܉UBm�_X��"������<���������@�J:$K!f 9^�{1q>c �L����,�D�s�_��trP���T@�Czz��3Gd��fX��֩��.Eܷ��2���h�LE�;�(?��Ņ;_�y���aE;#�M����=�A4ӧ!3e���0
P�@]K��$�[��f
�s?��ek
�?�i���K�2����a΢}^�K��ڦwaA��-�Cf/�z|s<���P��D �ICa���IF7K�܎�/!w�0H��#���>MUTzh5W�noKi̡]��ǗQ����k|3���;�{�a���A.pw�)�(s����ىP&�
B*K鶮�9����i�'ss��m�ZN�Y��E����ȶ7O�n���������3x����LE����� ��}�ŻxK: I��R��9���b�hJ���QxlzeE���Up�՟m�N00H�]Y��H��kd#f��?��u�u~|�����R ���rW9��m�7b5��D8�%EA�5��S5�%��!D'EK��D���<�Ɩ���J���-0 $�SE��S���?��Db9�Lc���b�	)wߘt�b�K 1��_�8��H�@�4��t��^����#����!���G��$�Z����>i,�W`f�?��?���$��
����3�V�9��������s�~٢E�� k��%H��k�z0����iS�P�B�E�/qc/A|0�$KN�+���3�ui_-�t�JfF�&-��u���A���D�Sx��2���p&
�]\O:����M�1M�Z�z�m�O�O�+�|�:��	z��%�1w��`)�Cߗ��=�pz�H_7��x�{�½z)�61�Ł��Z{����2q���T����3�[�
����%�x�S�X�;�˝��ļ��}��3R�+7�l-�_��BD?���WW;��q�Z�ER�xP�r��ι�Çʆ��-0~B�S\���Қ� $��r��Ǫ�JPV��I����ޑEY3g���bF)��=��#�F�	{��gǀ�5��S�6��e���˒�ES5|HH��Q�� 0̘ݾ~X�d�h��Hd�F@�t$ͼ����(�r����3�Fր+S�\�9>��?,������=>~�)������qE�Yni�r��8���ԾX3V��w<��[�J{��q�;QB�(�9589(-�}>�΋��6ɉ��J�-K���0�;"*2[��N�ξ@���S�f	"�4�?[璹��Oa�z�����Ϸޭ"�0@�}T��,%l��[��z��k{�u��g�F����� ��A��^��=λ#��+H�\�����9�H���ȹ
��N�,+0ǘ/�P�W&�A�#%|�_�{�h�"'z�幕(n����5=�[�%d���[�����X�Qu�2���v�H*e���uV�Ҧ,B:���:ܤ8.�wL
�7J�� ʟ_Qx��U@�(}�F��%'�W�a�h��k��⺪��������&�Y�� ŭ�ʢ�4�d`ϭ�1��7��}�sU�?ǚ_�?�ꚺ�|GU���sՂ�`������41�\jr� _�!EH���Œ����w�.яe�4eR���,˗�<��Y�y��r��v{�Ix�R{��U��Q��+��������}3��_���<�4]�O�K�Ϡ4��9����,����{\a��w0'٣����� �O������R��� �g F��w��Z�T�W�֮*7޼R�ɫ*���6x�f�V�����
W�]�Bp��wU,��e)+^T�����1��Q�oCr�Ƙ�UX:�-���:�Ճ@�B�R�t��^��#��=�c)2�����ξ�����4�I�_��s3ѱ͇�a��s��>[� �����$��g;��ؿ3��u5��8�1��&'�u�!��)��`��'�Nѣe�^�������U;�Z6�[�� �� `��e���*��h8���0s{_I�E�x���+ZH?Ӏ��}\e��<��`�3��h��Oq���V�3&���+l�t�J)�H|���AI|�'x��7��q-u8�l��5 ��i�л���Y�l��k}2}CA��X��3��[�:��R4�g�t��(29�_b~�������bV[Ӽ�'$?\��ՙwNc�:�9�?�q���%[C)������CtHɂ����i-
�����~�K��#�M�7*J�����5y�}����l�Wh6�#C�Z����l��y<q=d&�0�ʑ0�&���F�zv��Y�o:	�U|���Q�~iGK>�X�5V��p�{�"V�'�\�H�
��y��h+t�2��HYGENIhh[HI��9_@.OFy�lǤ����.n���LYu���´����u��G��TM0D�7��[��2vO{��MK��zW��KJF�˹��˂)j;�:�����D1����4�*����4T�uͰ����>�=#(��(��Dȴ��F7}쳴-�CTy7�c4@����)�T!����7{�DD6,@��g�s��Zka� l�dhA�lⵈ��`!��p����!��\�K�(��Oei�P����d0j1{���N�8��L:G�)w*�3rc掂�R���B�Y�����h�>�#T;�"�X�K�M{�2���ሪs�dڳ:��.�J��X>�P�|.��N3?����b��B�����X٨������V��j~�zD�4�!
�������ۇ���k2{��ly�$���sU��b��-���qk���G�OWT���:B"�2��j�!8�e���Ŭ�P�M�x��ڕ���t�͐<,�rZ�3/G�gm��/�4�X&��悎/a�����LL�!ϸ<�Q1S��F��yYI�d��uR@A�GBv��z.9��i�²� ^�ɧ��b*l׾c�蕊y�ԍ ?ey�4(g�!\>yųK���}���p�	>z���żL��ec�k}]C�dܮ��T���e�� $�w�������w)���y��^S	�Gd�=�� Ky��ơ��_v]�Rv�K�m�) Vʩڴ��A����<�ǝ��������=���۰�#���`��8��Y���%����\c1��g�p4S\]�&�Z��ӭ_]l�-�\���ry���T��sU�'�g��Q�u��~:Q,��PCc�+'o�X8p�\#��6o�in���� 3+rdRI`�R}�ϡL"�i3ew������H	\��C��o��1}�]��-�5�W�-<n��R��D ��9��5��tXw.�i�]g��N�]�8�5yژ9ƴ���
�����.��d:!v�O�$ �9ͪ/Q�� �|��^|1�<h婤F�s���xpLə�<�XōP�h��;��� ����If����h��W��JB�k�����WO�E?�!s�����D�t
/�y��l�m����6����&�V&�0շ4���D�Yݶ�l���kг�q��sǽY�X/^6��RҤs$L9,��[�,H0L�*&K��E�v؆}0�?���.Rћ�M�8,��?'���ni�[r�j�F�������)��5_�؏�<�w$ݝ����)���+��KJð�j%��Y���٩�-%�՞�������s�2_�Hi�æ�U~G�L�+%G�����i���� 	p�����#Lsy�8u8oӦU��굽U��d8��_E!�Z]��;uroA[6�.�A�����f�]D�u�&����p^	���,�������H9��!��9~�o�O~���=�l�.��