XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����9n�`e��p4�����I:1+�:���JI'P�s�0L��D����#�H�l/U|�o�6�t�=y�M�C�����R�0j�>w�<$&X1��e8�l/PP�R��΃�c���X�GU�(�Y��y����P��2�Y�)���N8|���6���+ H���H6��u�s�NӞ10ۭ�����T��&�'I���2���e�
s�y�X`8;�Y�m�)G�||��9ǩ�����6��7��e�7H9<�Zz*��D�A�#�P�ހy��Sf\&�HcM]\�4, �G���^E���N�3-��R	5y�ab�^���`4��CB��B��	��V�R�:μ;x0j)ak�CG�l�}[��5G�f����$M$tָN�-��,W��$�x��iX^���j�� ���+��˴[Hț�s�>�NP%f�Dԟ8m�|�`���Ml�n���������ĝ��-&G^X�A�v�ؒ].�b��1j,f19��i�+mQ��|e���+H�lp(������u��ދe�o����ۻS%������w}/��>brh4wn⩺����ٷ�>U�]�9���(��e3��`tI��,.�'^~hk9A���l4�h�^m͓уl[i�]F�R�E�f�q����<��#��DN� ��Í�$S�:�ڱ�oդ��1�K�dH����R��Qeb���/�;a�&�|��l��J۰�H��
��J9�Y6��C4�-�g���H?J��`�NXlxVHYEB    fa00    2040�����>g���ؽ��p��?�ST�h���<����z�\i����AVqpw��
� ���X�8����붍�sP2S�.Br7���Q�F��PON���%v�ڙ���I���������&��%QdD�f��O5&m�@a��VFD��T=�儈�)�4�0����N�w���W`Z�o�n�����d�v��/�&�����g��7�Z�:���?zF�J^�3��(@pt�5C�Gt���Ҍ��vZ��v��qGm>���D�Ɛ�b%��K*�Nȿ5�%�IFy�I'���9��!�����|�0�A��c�Ό[b4�_�����:��B�`1!!�����Y3hA(��iò!�_K�,��,�K�C�6@JA�%����s�n|]� |�X�b�ʧw���+��'�B �].D^���ubWYoGƦ߰�("ٷ�PLǻ�H���N�F�G�F����P�/ഒx&�d����m�����"�p��=��O)|�&�#��%wW!c� �;@�0�q�"ܙ�0��G���L�|�P:��y2���c�o
���g��!��Ůk����k^��O;/CLF��E
c[��B�Ž���Ѱ?�R��p5C*d;�����o�ܩ���k��V�ْ�z�K_�vQ�ѧp)Q�fJ�T��ܫ٫�l��8vI�6J�W3tE�)j���� j���/�6씸�]_��e[���1P��!�A )m�,��b�DA�`xT�ɦ?5�����U���޾J����FGT�|��dMbo������wzE��sJF�6����T!�F�ˑ�g&R���e��6�G.ץ��B� oT�<��/?��b]��Df��-�PO���-�C	ȟ�^;=�ǰJ�W���0G����� ZM8]����� =`�>���'~T��h�LK���M��Sfi1tK��x��2�ϧ2.�[����0+�>��S�����?z��qӲ�Rg���a?C��9�c7��;�zЦ,�����4�!��"�H)oD����庡�Ld��HDO#/�oJ@�װ�����?=Y�����ׄf4�u@S�>�q`7d�7jsq����?�gڴ_&I��a.X�R�Y ��S.��0�M�q��:�����v��WF_S��o�|,OBn6<��2�~eهbiq-���h�v$0f�ΨD��f��JJOIC�Z���h���
��p����n��g##��d�a<Cf�i��v���P�^le��RC���Wt7���Q����:; &�*KFiXj���\l�� �e�������r��n�8p�"�:eeK3-5�Ԁ��~�����8��� ��ޘ.s�Ev�33Jϴ�8O�����+�A�b~h>�\ D���o5��;f.0쳁�v���;C"J�@���]�%��>���/��<���O4�U���t���?�٤w��@�c�-c����_�=�eKeC���� .uAg��`F�4f�p�7"~%�֊Q�ʶ ą�]�<X���9�����w/�R��p�p�@C�<T_���*:_��YM[p WT�^�w����0�Y@�j-�*�E������O����Iv�g��(�C��$q��`���t+��!n�Vgɠm4!�$����"Ft�.��Ӟ�.�F.�+s�rL�0�ʩ�a�/�Ei�!븙բ,�c1��u�k�N+ː+%6��+��K���	�e�MgP��7*e��P9�㊪:TM�D���$�v�SSiY5$��"ySh��-�b��<��|�K��{�/ʀ���	!���]`U��}��G>ϐ���7�����ɇq�|��YU��
�������5?�h.M-D�s
�8Z���:F�
	�]�%��C��>%�\��	�O����R-��z����p~\�G�nt�7�E�]g�����(�<s���}�*�^2�[зM?�^8��WJ�&a�zR�\z��5���!�<H�����J�D�	�f��q�U������u��n���<J��-{U��q�"�����:�̖d����ǐ�Y�>�D���wd�		A���X����G�Q3�}D��x Dғ)
�F����f�ZM)����2�CtӅqk(i��W�B軽����J4���u�NN	D��S-@��t�z����^���9��DB��^��j����� 8M��PN�t&L���@!�G�&�l@0�Bc,�ǠS<v}V�k�I��LtC����S����N��褑�GL�Ky����"��;����
Nˈ=�� �<�����@��MN��c3����9p�0��j[��V�#����6���v��.k�ȯ���'����[���#�gG0��D:�嚂͓��s(�U�X�ų�̞����ͯ�< �P����=��V�Ø�v�����o�Q[���a�6���6��R_a@
�œp�L	
��W�i�ڧ��n>���i'���~	�z�Z��z�#2#�|V{�oU��Uu2�X7n8�$N�|�Oc�P���ۢ�y�v��>��R���IyLT�꤁b�,�`�V�j(���Cwl\E���RK�f�����䫄7��4��U0�5�Ғ�d��8́�Gn�#Xu?:h����2N���K�N�txоW�-��T�:��ߘ���4H_�����܈  �������3�D�lN�[�~&C���ἔt*�l�rd7�}2�������60O�-�c}.�;�ў��ɨ܂<��`�m�%�D�����1�V���28,�ox�d�uy lN�eR�u7E=й`u�LC��9���0�E��g\0���~@�7�M�c�$;v}Rcb��$\����>��xB����r��܎�iQ���D��E�NlEI_|��[��f�4:87�A�d$�?�LZ$��4I��䘷� ��d�� ��-�	����86�"Cy���.Y�#�@��:�p�ꏱ�ac3�j��v��y:m3�-2D�8;�$�y�b�8�ۡ�!جci��W�G-a<�r%9��'l�tޛ�"��5���HF Q�M~�ś�7/f���t+E27�\�.=� x>��(�%�*���G�����K�fH����u�*��]o�Uve

���0V��M�i20,bQ�1�}}�b:t��fN�B7�5z����9%�y���o�p�����M�;]�s}��Q ���Vo�AMx�Gz�tA/�:�i�T�ihTkLm��$����0^6C����y_��,����KWa�3�dK.�}������/��Î�<��V�b�Gx.ܮ�Cܰ�q�x���VU���z k'x���K�RD�.pvBD+�{�P*�d�+.��ب�uvV�V�&�l+`{�&��J�{Ԁ�j�삜j�^�H���~����n����i���e��fA'�|�Kv��W��
?��]@s���'ԣ3訳�ۂ�ݏ~C\�>U���� ��c'.���VYJ8�������$jiI��/����P���6�痎c5�ΐG��1����,E9�A��NR:�XB��65���n]�7���3@����E�<�.@���)A���0���2>��Z��y�6�c0������Z:�u����/��s��!P-8�����;��������1�-�e�E��0i+��n�H�[���Ƈn���3*.�C��X]+���I:DJ����\���Խ���1��+Y] ����&��F�gBC��{�Xv��Փ�}'����v����2^W���Ud"��wjێ��(��'e�Fi�����A����	I0��R$��BO��_���z*aoSiB7IH�������y�
�h�#;�Jh�.��aq�~�z�U+D^rt�_�[/��N9���㎛�%$�8~:QRR�P�h6�5�0��a�����W2݃v(�d�� ]S2��%+kq���Y��J'k)��v;/Y���Pep�����`�y�e��q�4��.�_�������i���J���B^�������s�)����f;�{��;�hE�䅟�U�� a)-� ��X8U��	�u�����rмSk����T@�Ё�
�;�;�g˙��4��I�� �7���:���E�t#���.�����
!�K�ԉ�I(m�ɂJRU��|�~��lȻGRb����V��4��]�����b&�Od�m�x�߆ʪ٭`/:mL�R�c�n�ߒ������Z�^ɬPBP����%(q�2�5���ݭ�/|5ԃ:Qo��5�����=e��m>���G�4�ܓ��Շl��@��b�Lx�@kidHˍ��To�Ӯ�o��-�/9UQ��@L�F=ax6�u��rC���ɺ&&��y<��!��-Wy���Q$ZÖ�7P4��ʗ�8<���Cr֢�5_���s>��_�:�?�  �RM ���7�]�]F�y��|ਡ&���@u��E/�	���#7�$ˀ���k�>�����v8ZRnY�|:��I ѵ��Avs9�j�Ld��1��
�;¬F�0��ԟ���}C�\T2�H:(p��cx��0J=�V�:ɮ���/�8��7�TB�P�#y���"����'��x��������M�
n�D����)��*H�������=��ڻ���gYf�K^WtU�/In������
��B
_}���鉄���ƚ�\�,�;�+	����2>�'Qk�d�.�,t�(w�2���`7�Ëp���������BM'A�D^�8�
�n� >1u�� �>�g8�Z)q��*j��H1��S�h�ὁBӽj�T�%�[f�3�|�I��\o~k&����. ��k5��b��=�r23�brEoN�}��f�������@$Ϣ�֖�DɂA��|��Lf��jФ��;
�����\�Ữ!�e�K8�p!v���������Jǩ֌�Of�~J�Yf�g]��k�Pk��$--�KF���0�(������YM\b�w��!�S��o��yx	T�ݷ�0SF�[Cۙ�PR>#���CU��K�))Pu<�,��p�PӦ�F���X��f�Ep�R{�IKhQ��%��)��
�����#b��5�S�P϶�rY�R̶�,$��;�٠^Y�xd!)��Z�[w���\`4�>h�5��l�mpM?t:6�&��-L��=��sVa���}ؓ�N*����T��X����,};��d��!P���y�6Â�&0Afϭ"���x�Wբ�_7c�fz��;�|����`��9p�Bv�<��'h��TOnj��U�֤�t[��J���CT���N�k�����Q�����,Ymn37���KT�LhC+.��`�A�~��5&<�B�eJ�o#s����92m����6�X�T�U��-7��l����a�7~	�R�r��Q��a�����=��� X�h�Ta�b�ݞX�+A���ef_���G�]2��:[K�Ιh9�u
�����(Zf7!Vc'.���D2y��o��� �%���NGu���r��"�V���=}�s��^��i��d� l�w��,���������[�|�;��$��~�O%�,������R;|�폈�"�Ч�W�%��B`Cj%w�77���~lƂ�7��l�ņ����jiR��_R%Lڪ������wp��H~�3,M6p$]���컹���?*�N�V R�p�$ی�:�F��������d�l"Tr�N"�`^�cw�1%�R�����B�d��:�6/Qz3�!�]*qX4u)
^ �J���\��)�-K��m�+�cgU%�vrC��������t�f��OΜ���9T;���=�[5����#\�w���zv���z�����+��ț�V4,I�d�o���R����n�ۧ��X�X3����t�δ)��D��7T aO��S��&*akd)���_j���q4���Qo���n�Г}ઢ�"$��Q�ԉ�# ����Qw����#�ۆ�-a%8��GѡX��R���s�fpwV��(�Ed��W��L'}��;i~4�;�f���fXF0�f��C�����(�ڤ=I&#�O��Jy�C�W0-���i����@�{ߠ/i��9�y�=mI�w��3�jTPd5��v���*q%�(8�h7MwlZ9��F�:IÎ�	���U6��=Ђ<Gh�j����.$����v���ٛ�����h�'���A�7��{胼;X�����"I�aw>u��=b͞��W/m`N�U�6��$�֜F.�FtE�����xe	7{F^S�!�_0�(�#�5��U�4�h��[��O�/�;d'�%N��#�X�`�UF��h[Ԣ�+vg�O��&3:�t�ѹCӬ���8c�� ��5&oY��4� �z ��k�"9�y�p%�أ��~$M��㛡w���qY Y��K2Ċy䍟b=P�Vnq�t�L$����bv�o�vG�b��\�gba�N�2x�㳋o�͜���]aX��{���u�b��ae�G4Ą=D�8S�Qs�r����ѻU'���vQ��I�9n�8�/Ͱ� �ۜ|ُf#�_���v`[UUw�s�!v����xS �����G?ݘ�+JJ��N�e���C�����$uWr�o��F�4#j�"���i�
�֮��L$�!�y������Lg'm>h3Y�I?���cЉgdg20�zU�`��m�bSjn�
A������>O���}�+<�㔯T� ��9y�flK�8ЋN�S��(��VQJ���IK��(���Sm���ڬ�&����}J�<�a��3�&H	懋���sFyU?�SH��ч+�ڸs������#����C[�$o��M��L�t�y?ĥ�ed�Ū�����l�K�i�1��:�����
�9�x�A�qm�HԨFrb�+uB[���so&�:�2�oUk�NM]�j6RV��\���D���̮����.�:�wݗۉi�'�c��~�*�n�{̓����~(nݓ�sy_�&R�*k�X�}Ta��z�d��Ô\��5�NM�:�<ޕj�p�H��tɁ�s��CS��ò��N[�iNt&[l�+Uk�����h�ը�t�:��)����˪�_������\���.Be� ǘ�����A�N�,����M�D��H���CgfѺ�r�)�y��孰ea��K��{��e��)fqc��2_�iۦ�2�������C&����$;���Ѯ5�(s$i��"�%�w%�Xy�ϰ�7M�ڻ��%�&�˷�lP��.6�tg�z'��.z�ط���Ad��R6�!�����q����.� �e�'�N{�F��vJ[�]7f���ҩ�AᲫ��\4�$��+�Y���%@��N�Sck�$��ݛu)Ӱ���/L�㊜��/�lӯ[�nMU��I�8�5�U4�IL�;E�n��c��(b�#l40�LŤ݅��}dۗ��������F����T�8�|b�%�NlŠ�_l��#p�V�?8��Ԉ�6QBk���)mn<�'/�Ń�w,ɷK���q���n�B �z&N�Io7��((�;�
���ޠ���?�{��X �TXlS���������)C�94努Z����@3'ϸ���eڪ8	��˙L��`��� �	i�5z �"�&O���68�Jr☝\�{'G�+�F�*���3��y�#W��-�e���߇����%{�bX)�7-OL屗����n�ࡇ��B������Q�R:��+R��eV�����ĵ.����5�-�U��q<>7l��!���M��Y�:�Y^;�H8f��	����Hi��"rb,�y�9�ș\hAc(/�mJڼ��_T���*3}�&��{���5oj�@c�zr��sĢ��bcW�*��`3����d�-��ѷOp�]����R�A��n������ޭ�w�����B\�ka�P㣵�� ㈈w��Y��*x�����o�����a<��*��÷��MD`l����;8 gC�)'�-�7���Ju����;�C|��=p
D��}?�!q�ք)?9a�$t�	��M
�2%��78��>���D�=�7R;*Q<�@���gd`�Yl����;�b���3����ҩa�+�\#s��)���XlxVHYEB    4f62     b50A�m:��Ҕ�VX�d�R0:�zU�[�$T�y���E�9��s��L>�}��$4��4�@;�7�Z�Y�_�G��آ�b���nH/Ds��n^�~i��$�ww�e'�weWH)��`�9LU�C@��e�|z��I"v8z$�Dtpyi>�Z�r(y��}K<�FϏ�(�zs$���fr�)u6��G2B�XWB?߉q�˶k�ʗ�`�6�\$��'"�\U�t�.����S�rɐ�M�?<����/ծ��"�#O�И���P>���)�y��Q0����o�w�LX^�/mr��ۮ�Ic�+g+7�Zbh`���Oo�1��_��B�*�iw���N��$d2V���ԫn@F�>�y@93�����Qq�jc�����_c%d�!������xZ���t�?�����z�վ���޺��"�����O2�ڊ��`���w�˘�caæ��խ�
v�~ۖ6֔VeO�Q�aAP=�)7�嫀/��k]�*R�,x�>����CJ٫�E7�L��Sp��<�
g����_��j��C�C�Q`FL��"R��Ri!�����b�e}-(�T�m���!T�K[!�~ �Q��� ᧁ�M�;��,�`��D%��	���4��l&����@��#P���rT��T-��� 8�D�9����ʬ���f] ��.&d�x���:l����=u~b��q� �:Rp���U2�pد�>�:�/�Wbc��R�ka������������������Yj.̚P }<Z0����U6=Ҏ�L�n�TĠ�sK�,�3���e��t��2����v/�n��ޫH�;��ڂ�VH� c�Ҝ�[��u`�>�-{+H?�__T����.|�㯀*KAPDr���hT��7�)���R%'��R��0�q��X"&i���y��>�[#�w0O����A��[�C[?'~��ܗL���͞���&l�s�:;�-B�Z?x�?E��;U�'��ʝB����'�Yg�0O.Ȃ�Ţ֢�Ʒx�+C$%�|����/���c�=@N���U��Z~�!TK�{	JO����-�ˉO+%���(��<z��Q�E)rLD����4���F�q�k�-�������L�-q��N��!�e��点0&~�g���g�Bc�&��M����S���SKRw�K�K�#Th��n�qR�x��x�H�2���!��M�����3db�Օ@laKFHa�����i-�����D �#Er���`k�:b�dhN���F�Q�������L Upi��"�7Nd
g"?���37����'$x�vN����y�z���d
�����X6|�K�%7��H.	
����C��|}Q�]u��U�o_ew)��:LV޾>���O���j�]ͷ]-�G�����e�0Q����2���m�>;��c�y�)өbS*敁�]�ۉ��`ɴ���-��;�2g;� Zc)l%m4Λ���$/�%k���߿��a�6�<���ϠiF�X��o���fٚP8uo��:��9�Zx}�e�,[;�M+��%mD�Zshm�����f�C��ѓ��R�6��l�k1�y@����{�����oV�bbaG�R�?�-�#�B��J���3ƧW8�c�#���ؚ���\��#�
�� �xP��z�l^�E���t��a�Q��l�G��jK����ÌE�tw[�̈��Ɏj<���>�w%��8/y�B��s�ܵKcL��qZ��6�s�T' M���5��~��R�ɤо�z�M�'�qAl��D=՘w��s
S�����\�$P���n��Ǭm?�oꛈ�ZP '3!��0�X\7*�HnL
���0�7��{��o'n�cC*U�H�w�Ր2>����S�k�-�^]]�
�����O���FOo�ӏ�NyC��7&��O��|���5�%�4;Vς���0*I����1��K�7;��sRQ{1�M���2�% ��
�6H���
�0;k<�U�Ul,vl��B伂ֵ�n�^�z1�"Uuh>8Њ�+����_��9���pe2��ֻ���Bs���32g��W�9�ڴ��m8�p�=��J��+�UBr1���3��f�
�j�/@Mx׉�H.����)I̾���,}c��O8J�f����w[i'x�7��MO�Q�T� ��(��5�72�8���i�*qEj�����*��U���V=�r@+�J��x4,�|�l:���a���dL���䊎���62T�v�Z`[�+�*�m��~��k�s�g�t)��. 0y{��yCI]H0ɸ��rl���"e�����S|����؏4�:[���Y�=�r`�,���{�tYf�	ї�ê�}%�4��(�88c׬�pf�\=��/_��e����1'���z���Ϳ�V���T�7�4��V�O�� ��]Z�v�c`��o�;?�8�&�h�+��
A��/U;��Ӛ��K�������#s�L�*��@���qh:)Pq\������]lc��r��I�lْ0F�F��k�;m>�21_5v��m�.K��r�����;���E�jC�ԘHS��	dbUw�ѤH���`$���,Lù��v?>=�nX�+� ���n|�T�`�v�_�G��"ν��<D�Q�����$Ѧ���$�6ya� A�b��FM���������w�p	�u_�����������L�& $��	�Ǥ���U���p76�������rΞ�C�����U�"��f���Go��r�\D��G�O�q��g/��vB6߅6/�ş�`U>:�m�׫E��n�rf)�}>,6��+�2�?�