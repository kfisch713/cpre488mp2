XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͏8��W�	qܴ�u��VRu�����&�9p��Mlc��{�T*tv�'q2�7���[p���s�賢d�R��[�]�}��t>�ٜ����}ئs��3sR�܈��2�N���R
,Է���I��#;H��j�j�;d%�M�ܿ��74\�ǎ�",��*('�<;A;pek�`v�D�#�j�!3̭͇;f�Y3��Ԛ�JEE\��c�(�����V�,K#�+:���E����f�,Ȏɧ�f��A�*�]������u�'�� ���c�����a��:R^��}�(�_��T�^Ѕ����|�bFO�`��+�	s:#����X���]
�a���jm�)F+ #6I��Ĥ�A��06���/'OҮ��h̡A������+���K1���b��:bB���]���e����@R|��Z:�v�b�hfy�X:U�>4�8�D�������d�y@��;�C�u�mnS��-�'� ��DV4ĩ� �y�c��V����� 3 �K{3&�_��WVZ���D)|o����z�m>�ʦH�c���8|#P�t�}�K��p!|�I�k>Vu�#������4��=!i��0�����P!��	�?�j���L*�U��`6�����j����4,�����2t�\3�#>��AN$ߊ��u��`6<���1>�.,�� s������Ibx6� ͘F�8u���Q�%��5;�Zp���u�ir�y.h���9Q{�!RX29ٕG;�R߫yf�w��փ�U��|)�7�v��XlxVHYEB    2326     980�}�N�%	D*��O���m9L�o�U���^�Z9+��9WY!�2Mb=���D��=�T"����������8� �g>3��w����񖯡e�����wԴJ����%9����]#HC9q|��,��:�����y}�S��� �\7��+K�oI���%D�.S��Ӆ��_����s����a����~��h#A�r쐗
̗o��È��[F!��~�9��桯˥��{�T+��}u����#��h�t�E��p����!i,�j���/�4���_��Ny��6*X/���e�I��X%�t�9eV4M�\{Y�.�G��S����� q>rĐJ��Y\��F�����F���GW��:�Cvd�����(ۉ�e	�[!t�V8�+`N/%	Β�k��l�V��;`P�$
.L��@� ;/sn���.�TE=�4��B�>_��n�dX���t	�~)J��0����6��Ng��&�b�cN�F���9�Bԙ��k=5p���G mx��%~R��%��)<�D\DC�N�!��cn�	������ L+�s�!Z%��u����*Tt�������rȡF���Y��&��n�noU�΂��?��l��1*�ܭ}�*
�[{��ю
By�#b����#nfr��]tl�8��LQ����sB����AX�ĉ�ie?k�[6�)�o7C:{��K��wQE.���HP��Ϣ���T�J�I�yy�R�H��B���05����G����Z��鲘���>�o{ơ���#$���}Ǉl�S8a���N\���0��zz?Y��������ܴ;�sml���� z�`���F�|̳9���Ux�ފ]>r��l�6yS������-q~��5!��� �e����<+�ּ��[r����Q��>me����t��O'0�EY?�c���E��{h�x���q�b�$��\�����oŌ����~�����VJ'��. �#�S�O�%�4N;h:�G��������z����Xq*{�ؤ���%	|��~u@�@�I���6�l��h�0Q-r͞e�Ҭ�W�"3���)\U��U&.�F����[�q��M�C���S��l�M$G�)����?(�*��������s��j�w0��A*�E_@�n��0��ƣ a0�At~Z���E�uӕp��m�؝�d���(����x����R�g(���$�ǲ?�#�W���C&e!��r����������@��?
��#up2*�w5Pk��d�k���2��=c��p�g�gP�s��;�+���Q���e��
.!�Ob�ah3ڮ��d��1lI��%V��1lÔa#J���Ô���b��%��<Q3mM>3�'�vk�,��l�V#�ԆT�?S Л�U��>\W�g%��)����4[V�>Y���j
����{I��Pտ[5e�n��UI�_�zU���.,Pgz����佞�|�B�L�Ti�e�Aޑ??���ǲ�QqY�7q�N�*~�kp��9|e�����'�|�>�NM\�vV\"`�{l�7uٷw��w�����u���|��Bo�����(�:1��+Y�Y������m6�z���>Т�����ez����۔�^Z��_1��K�@�+%+�G/�̰�a��a����¿�)XP���Yܐ��Ժ���|Q�,e���W��qY�͕��o�.%��$|�O{	Ă;�0N�2=L�����B�4�N�T����Q�	�1"��SF�8���8P[�v��2iz���B4�݋��j�גE���1�u�9�(�	�)?��Re�H�N��4�C'h��P��}����HU-�ĺ�ۿ@�ږ��X�?8R�D¹�Al1�.���?ÙeZ��jמ\��A�:��?����n_������9��ש�6����q�w�[5)����!����Q�8�o�P4`d@y�l���b��z������x�h��˹^svck�H":�u���sh&P>"�+�נ�m%�C^��8�.�!��ҿKD�6f���>^� z`���:�nTi�n�T@g�P�܎;8/ܭ�������5���P�&�C��BÙ���l�l�CR���|5"))4�D�m:lӟ�eE�A!-�V�s'	�D����#�Z 6	���L	�$���|��Pϼ�f��u�M����}H�}�]�b�"�+�!­b��	����c{�g��؃P��>���ټp��ϋ�����1����]@�3w��drgJ>e����`	w�r�Q�?>3P���A� ���S���@���5�TC�W��n/ld\z۔��E�X�S�j&1�;�L'�9��5�12)�c����-0Ĉ���!���GQJ`�0���UQ
d:�M�?�8����F���$�����Z;����}�<`�&�S���:D���'�Fq=�