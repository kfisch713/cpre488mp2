XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��em��Z�۫��/͉c�N{p�.�P��;��ދD���ch�m��B�y�3ǌ>3Q��#0I8٧ ����Ezw�֮װ]��B��H��W5^q��(�d��YHP���#x�����IoU��d6Rpu����[���B2w��RtrԈ�w��7nEdQ�Y� ��^u�QIg��;�K��P?h����8O�0|i8@�X���ˊ��4R���!��$�7�t�j�F�R���Q�%ca٣�7B٭����jſ��w=����>?�p]i��M0!n\��~sqVӃgM�!���;s�n>���U⮧��҃�*!!��l#��h�\��i��lۭ��l�:8i���cC��N��
ś�FQ\�+����L��uߚ]���X}���t�$�d�e�|Qa��Lh"�@̚�t�q������d6	������6���	>�y
c3w_�T�`�m�g�vd�#JԲ̧,�ev��N�*j�#�ɲ��$ף��؉B�(����� 2p'�MW�ֲً���w�0^�|=�ݭ����@�WW��/ā��R���`$5�u�c����I����iQ�Pe '��%���j
|�h�R��>��OQ>(���jzQ��[
\&ɧQ����Vt,�J���_ɸ]p��o~��U|���ĭ>�T�<�܈�4M~/*�5X��I&�������}�mb:�Տ���d�Q�fI�lu�KʄF�E����J��;t(�� ]��JK9�T���b���?ݼ���\XlxVHYEB    2b75     cd0N�T��_	��ȧ)��R�����%�,Z����(na�{j�"2�P"���t�8�٣KG��'�Z��bN̀@��C�~�u*�M��x,d��(�6��}Ŭ�bx�0Ѽ�����̝-����~��ى^1��j��q!h�4�69��Dj�`�k:��B�����|	~�g6�x��,�@	�Qe��e� ٲ~�K�(,�V��m!�s��Ka�BbZLW6 \M��r�d���%���'�Z�h��	�"�t[��-��;[1I���@oj�e��73��+Kh�4܏�"��~q�
�� �ޚْj�\�`�gVk�P$B���y�)��S�������/�Q���Jд>�����p��o5�چ�}�U:ZCT�~=�O��A/�^�fHz�%��h�P��a�������d��Z��]�cG�����7]N�2�ʵ�!E�����;��D�J����Q����(�ySt��)��0|�������.�y�v���)7V��T���S��3'p���^F+j��}��x�� k�b��]zOT�"�g �0��;&_8gj�(n��绬����+���z�va�@P�4���c�룞U�m�_g����>�c��\>����ɊK�A~)h�,�N�A��)�h��Nn�r�hh{
g{�e�R���\�I��[�\Ì¸��A�ʓ��W���
͐�g���a��ŋ��I��c���.��x�P�&��QH��2�+��7VUy�J��5a��Jr�}=����]������Fi��G���oy҇DV���ت����ٛ�cL"�VF@N��PH��]�3��x�����1�5��/*8Ҭ,��λ%Fay$������"�v&6Ēށ�����j$��3�4�D`S������,�/|��y���+��C�LѬ'!��tu�'�LtB�5ʄÓ^6T�O_1��5[�Ц��P;�|W��YI3���8��.�H�HҴu��TEӎ�uE�tl���&�έZ���h�,�+��i�Qa\L4�,���?ԁ��21\��h ��=���(IN����&D@�l>��%-��,Z�.���cF�N��
�ct�ݷ9z�B�u�罝AKvV+9�2U�nr5j�)5���EK#P\��ykMT*q����ХpI>]w/����}~bTF��#��CM>]x�~wՇ��]�?J���ψY��3� CD]��b��|_��	p��K���&tOr����I��3��(j��!
t���oGH��"��2r:9�9���4eY�"��AB5	L��ҡ�⊝�x�ɞ�"�Mͭȷ��:T$�� aU.�@i�g %��u�n����=}Fh��%Q�
��*K���aJ���T�i�+wvZA1I7��� a!�lS�P�ʖ�=>�Al)ԑ�|�ui�6�^A(t\�z�
82�C��� �k=�'�K_����1�/�{��QEb�E,�h�;�9	�$o�_�U���8G���d-��(�B��)sm�����@oź�v�@0�G���p&�!|���#��cl��=�m����G��%E8�3�v��9/���ȁ�Z%,�`�gb�՝�x#��w>+�H���c�;$?i�`|N_6z� ��<��Z���{�9h�	�p#(�[��Jз��-�38T���d��{K�Z��R����ܗ�g�x�N�MK�tN��&��4��rx6���zT~9�g� ���@ĭV�%~aN<dW>L�F���"�Υ�˱0P�3�� �I�� p!��p� gfԹ&�!9N�����G��f'���:c(>�k�fÞM|π�%́v%�Q��iW��"d~lHa��?��aA�{E/?��),�T
���v�H��_�n%�V*Hl�U˪I�����YHlHs�a��bF���CؾA���M
K����$%��\�y�~��TWb��%�/�tz��狙���	��� ������)e/$�z�g� �;����h�hÅL�DO��x��|�g�e��ȫ�M~���?��EO3d �.�u`+4$�����p������+
��+o	l�W�������܍���}������{x|����P[U����� �6��+)�H�5�� �{5�~|��Q3_�s�����O=&,���7���Q��5�I����Y}�*�@�I� ��3�)t�e�o?�Kۡ֗q�!55�����Gx/%c&Z�U�����J��|3������?��IE���C�gЃ�uE������Z���A߻����v����R}��J۩��ϵj�Wf�oQG��dR&�XB&��:�)RɌm4OV���4�s�t���{J����Ϋ�W��-WVMg���0)�暛	o����� .�3������V���#rǱ<$-l��  ��ٿ[�8�J�v��J&��c@��������� ;��8�G�#u�pz�20�<�W,4�sH���S���I4o�l����y����%�:)���'?>�=#�룾��1�I����`�\����Fƍ�B��'4�wq��ѝ$�c}��So�RN���h��|�g��!�94���s
��R5����!�b�֟��3��yK�^\����<WkO��Z5��'�K�	���ۍƽ���n(�e�+�zt:�=5;H�Xx��ΐ���V.ߩ3mf�M�.�%���K���ia�PB}�^
�������v�Fj*�Wok�0���"�VZ��H���F����� �R�~�W��O���DfX�7�r˘J�%�/>Ћ��ê��o��-11�Ż5˲�fg���$�-�}W�
b�%���o2<�IgKf�Y3�����z!�!���o kb"��U�ٱ��1�P�3�%rS�K�|f�8�Ubʽ��7�� ��X�����A�0S�`�y-��4�Xoo����~w�f���j�ߛ.�n?:�?9/q���%�$��G_�������ƕ���cEfH��� M�O4��=y��[�J*ӎ`b�Tv���!6E������F�0���4��hdOm��ٚZ2���{3�'�I��E�L�B��2Y����@�o�X�g9w��&|n�����H�%x����4�e����G	��Ҝ*���.��a�I�+)�	�Ś�Ѩ4��z�~����]����j��'��ɝ~�VFi6������y��j����";!�p��Ҳ�B+YȦK�@p9�&m��p��8!0���'|��I�~A1���