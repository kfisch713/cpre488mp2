XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&����G�aLA���la/j�3������)ak�Ŀ�����Z޻?��	�;O��J\�w9�����9��+Zv������9)vL��\�,ӅU83�>2<*�8ݾ�#/� G�g�cZg�\�����ڦ-�4g���=|W+5�ׯ�O�ik l�G�U�����&�M��ט>�:b)�\\��I-�C�k ^�|����IXw�tZ���
.r��q5��+�ń�`�=�X����+@��ԉ�8Ƒ)r\��z��f�P2�Œ��d-�A�����1�^��g����L0E�b��%�{���jzr�=���CH��Et��߰�\��/�z�`d�i#�v�2��c���3JK���zۭ�`�H-��p��jQL����T�P��f���v$[,����)XP��|�]�9R��s�qpX7/�zi�:��O�'P�
��.ٌ2D��C�7_�j���\�m�4���%|�H��t�F�u���ˇ<fٲ����U/����,E�h,8�w��+���W�ؽ@OBʥ-9J��������!�(���G_�*�M�˓�ε�����^4��ɩye��l{!�n}�}�ˣ�.�r>��'�Z]G��m���dt����j����,����d&	�Jc��Š]���c�c* �;����8�2��Hz�x�f	F���Kb�>b��:oJ������$c����k���F8���Wb�P��|����"q����PLc'�0�@*|l�A�f����-;�n�GHRa&D�XlxVHYEB    5fea    1830x�S��U��Y~�d	kg�Տ�i唡����f�L���&�����
(�m��V1k�L�#�
~	Ð\��],oṁ�7����9ϝ(=�'c���of�0U{`���]�����W �%D�DЈ��,�Am���gPu/�5�QJ
 �Ȼ�����Y��$+9�cA�{��T� �_�@4�+A
�<�D��yq��ղ!h����G��3�[�@4++��h���8?�YT�{#�o��֮HoV���[�T�hl�%T������ꌵ�X �W���Q��)[���q�]��%�B��h<��D�u/��A�H��v�2�nZ���p�������G��#.�lO���e ����c��p��V%�<h�E>hB�!9�?�<|Đ^�)����7|r�w^|��K�O��uhpw=���CƍӼ!���yl=�.�+hy��:\#���pV&����x��tVh�����
S�������s����"���SG��n>�w�(�῔;�{U���}�0'5����E��P��<�
�G��%jS�����D�=N����k���3u�E�,�"�i-�!�;)�}ż�W��3k�U��z��f`د�b�ض�Y�-�sVlvt������$9A5x9� ^������_qN'8�4�
R��U�];�(�X>m]��bir}0����F��0qJ���I����wz���k>�ݟP�Q��R�����Ǭ�Sל�Q��Aęp�u�\�����Z�ܒLٲ�x1"��#?��ܼ!y��遛�}��'M@��=��]ʂ�7�Z�+�=h������Qz��)8��qA�Q�#�Ix/2�Hٱ�o�S T��q��z�(�/������*�Rp���&� �o7�M�f�l�+��e��AE!���%\q�Fd_���hA���&MBt�	�~Bևp'��|v�Hi2Psd�Ҿ�rjwMFJ[�4���Q ~or���:�S��2� �t� ��;�0u͌��٘&��I؂����[���~P�~!B��;�D;�26��u��<R%�M�� �zA&������duk�!�i����M$��f�K��8�!�2M˼*��*��Y=ࢯ^)�;p��e)Nf֊��g�k����l�qᖿ�~Vj�p���Z6?�����[HqՉ��3�������L	������6	6�u�0]O���WY��Б�ӱ�C�f�LF��w����7�J��V��=������'`��E�Y�Jl�i]߳!�P�7�b�����A|��F㱱�Crݪ��Y_��Qo.�	�{�3���p�28��a(n�a�0<�GDq�D?v�㴽JT��L��T	}L���q�-n..��ORo���u8�In����:�����4�xu��G�Gҟ�~��za-�w�E��N���}���W�pT�b��B~,�~ߒ�+',�v��.t�v-�����`��8�WZ$%Q�C�!�㟊j���\睽��_��)��	37[�g�k����b���{H*�:ܘA1���{Pf#���L!�y_^�TO�!��/Q�+�#��s\]͈���{�kF�")�ћO價k�̶��>�FV&�%�[�}�YQ�\��'���Wf��8����I��';�Q� i��>\1�.u��c}�ARA�+��#�ArQP"���\3��_k�O�5���c�k�<~މ���$5�Z�񣱀�0�9X��3b���[��n��v�.����泺N��w�Oţ�g-��v�H������R���/v͗���E�)S�H{�f�a+�rE4,\�K��9��|em��8������W?5&k��&�Qo��0�x�f �zｵ����Y*s�+O�Q�B����]��?1uR�d�~�XRT�m6��OـFqӆ���|��X�}Y��]�[2\?�7� ��3Oi 5U"\����CN~$�eX�ԯ�@���qf�e�Ř��> w��$+D�(z�����f���1�MVA3��q�]�-��ן��2O����`5iej�*���]V���*x��W��c�T:CAz�2�ڷҚ�&6�o�A�0j����O>c_����(�Z�� ;�M܇�� BQH�sj�ϊ���B�:��iD��3��س�}��!3����:*_S-c*8� �~���Y�	��д^)��0��w"Q�pth�j�C3'G!<Kvm��]P8�%3���`�&�@��Q��g�zHq��f����	�w;W�P�i�����>���Ǔ`R�j4G��ǟI}ojw��7;ӳ
h�]�*`-aL(5j�RYOj��6�U<U�l� � �!w(}��Ӣ�6s���	G��&�5I�Bk$^�^���"}�ͯ�0���@kO������+H�E�n(	�Y�!
��|���6eh1Έ!��(��h�(����Ei�K��P"8�M�WF�hr]v��p�o�9T���([�G%���K[�ؽ���T��p<k_����k��O�	��k5�.pܿy>����0��n��ǟ�r�Z�cZ��g�+/GC�d"���NR?$�9�#c����g�1��2�7�����6����x�`ŉH��h'_��~�a��8�Np7�Fh��Lަ!=v��b���dR } ��S=]z�j��y���I�W}̮��gV�iz�%��;?¨��~���	$�1�mW0�Ú�r�e��+&w����U���	��!���i�{ +�3��ٻ���-��#��O@�[�7p�k�Z�re��ǅӔȀ���Ok/;��ÿ�+���dqDx<Nj�P��dvk�RL�f����C���j������P��ּ&���e���
�7�y@- t�_?s���3��@����>����XZ��L�˖,��r�߱cQ۬e�m9��Z���\�$�2��_�!�u5?�!l;��A����Q�)z�n�92��į�����0JV7+P��KV��\���.i�b��Y�b>䀾'B~	�Ǔ�{� ���a��?���p]���f_O�(��:���v��,�ۻ� xn��t��}^w�>Zȕ�²���&4sDoc6�q����B%���Wc��vyo�R��#U|`_=O"N	'��8O��s�����a�z�����qJ�����Q�����'�T�����N6$
J�j�5=z��^�4��R�{/����2o��c�'�Z"���A����`�<`�0�ؒ�@0p�5/sHC�x���V���g�gr���4���� T�JٴՀG�'���\�U�3��ל9?G+U�Jifٮ�9�"M��Tǽ
7u��Sމ!�:�˦�T�(&����0|��2�n8tكT;5w�ic�R�_k�E�$� +ë�јҠ�"��Hֿ��7T論rVO�ׅM(���#l,����*�[CJ9�Z$�y$�I�:�i�����f�A
d�I���h�AQR��E�����)pM�����n"�j��#ٖ�����$+���>�L�
��)}Y���~�}����݇ly'��ln
K����|с�a��2t'�#*��Ѱ&���ģZ��O�q��N���2êCCS���Ļjk9��E%;��i�/��#�h��y0|���Ƌ��k��t#%������
�!�M�I���@��C�_�U&��By�Ƙ��4�o���7�c͞�����`y�����$ū���]��F�v�ƙ[��h�h�3����7h�����ٶ�S���XE���s|j"bq[�O#�[�,sc>��Ԭ���"ɉr����}��������"�/a6~�>*D紛�U���,���MV��7�i���CZ*�NNC�i�, �ӡ��k���F�[C+���o&M���M�W&�Ժ����b�x-�TS���~B�W�C�h��GO�VZ��l?Xoێ�Z��
��C�n��&��B�8�k���o���)*�n�����`m��ݑ'(�Lа.�9N>�:R�B�_���>�̈�q�-�"�^u��RW>�/�mXw.Z��:�|��e~�{�����@��,��h7�j�QC��Ȇv�%U���I8�R��yH�vr�J|(5�<DI:�g��C��|�࿈\��I
E���N�7�⪄�4��ȘM�!��k���
()��[3p�zt�-��8-���]�@�h`�I5����/P�Qxm�޶&1�}n�lƮ��w��0R�x��=f�!K�S�ߝ3��������VŖ�I>�t'��|�e��������C�D֔#�"˟���&���vM��o ��L�iV+�,|��n�Y[�.�qއ�	��OY�A�fhϥ>�"ɫ���iʓ] ]��4(D�P�M�a�n�u("-��prIu��0H�!"�k��1���݋��u��b�趫3p�@�@�� �!�j�q�)�w��s��$ʙC0���0ma�YрUc�e7�+�o9!�i:}���K�z8Kq-�k8�z����{�d���z��)�.B��a���_	#f�o "���T�mhooIR��E�AhN.�z�俺/�|eiN�$$`�C��7������G?tW��)bᭉ��w�5cu��q�Ve������h�啊�HIjI�^,8�~%I�q!�L�^i!R�R�t��?���æ{ȑg+������	�ѢQ��:�����&��f�/"������+�
���0IL����]��w'�6]��)�}7���	�����w���>��#6�����y��A�{D>�IL���-����N�h^"��,���K�@��^�o���B|������a�ɐ����~�d�s��#W��H�"͛'�ǐ�N�3�yc�
L�������6�˗����b�zu�������/I�Iuz�����.U����8C�0�f�.�1�"ʟy~�ڍ�-KePk{d�6{a�sg��gu%�ecƠ~jw�d��9�a��t̆b?�6l�"�k��"5������x���P�B3A ������\氬��������/�O�w�݁y��F�=k�%	�>��w'��at�6l@���V9�AD�&��|!���/R� �yW�� �#�N3������=%�1$qo��6�	�భ��2�ɇ~������	��\�e�{*����DM�@J�A۰�y�;���į�A�l�Ix���eE;$��KL�Ug�f�QG岏�����Ԧ�~��]1���h�xϥG7�,�(�('�dݬ���� ����#:,�u�̒/�����v�I|�,��(�m���A\��c2�=���O�e<�������|�<}�FF
[�#N9����}�W��c�{6i��2�  W�c[wb����+>#�s��`���ĦsjWG�`_ӯ��aqzc�>tV!�-G��j����N���JM_*{����
%YK����Z�
P���zv����H�ùC��M���:�>���`��=�ˌ��ʠ�zA���xlel�� [�Sq��R��1��"�F�`�Nԣz�L��	]֯s �x�����Z2�@d+FWH���������)�^�ԣ����ҟ5�H;S��T B#�������y����F¹����%�\iǘXd����)�v���9��?0�/B�$>�U�M�����D��"�4�扯�,Fa��j�/�A�#2\=1�7�іnA��E�Sz�ʟ��*fh@�$����@�;z����m~x�M#�{�Z�<�1(�X��|��_��{�{���Ԗ:���FMڃŕ��sHot_��_+E����RJ,kAL,D���u�;�I��N�gi{��1B���X.p�v!��e-��09S�V�Z膲�B���Ɲ|<;6v �6�����͔�c�&3��Q���˴t���2f�y�c)P�ŻJ���ٵ�(�X�f����oh�
�'`�?��ev���OJ�A�?�AJ��/�Q�O�A�8�]��Ƙ�v��U���_ǃ�ARF���oPq��0�L�U$^֗Enq^�v�c�)W�}l�����;����x���F�=xL�����E
���5����c���B��� ��ݺ�E�_o4[<�b��Έ����N>��D*p
�������0 �Z](�ꕄ���kч6�@3l��' 4D��&�ӄ