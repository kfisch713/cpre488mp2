XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������l2��r<c���C?�03a��J��&N[	Ϙ�a�x�˘-k${�r�&Xѕq�2�X^�r���Ot��6H>��8�@Q>����.��_��D:�`��|wзAr����J�|� u��@�3�ջ��]�.�z��{�L��#
����mAT��� �2�B��1$q���.�D�?Y
�~g�N�\�^�C�}�xd���6�;���|��Y�3��L�w+OiB���&h�m��ш�^��rzQ}2I�ϨG�,����ɗ����,��/��&�N�b�}	ڵ�DI&��]�<���	d��t�*�g��V$A�_��G&��}nad��@|-ss�ǰlYoH,C�W�}��y�jT! ]��Z�L/�����O�ke�nu�_*��Ze���Qլ[��i1-���.������F�!��vWhF�o��!���e:(�1(�_!���3�6@*7�/XZly�_0��TNrd���^�f|c��X�<@�>�E�\ÑhWr7� �!�o�8�XH��R����J����� �&�\)�@~��MB�^�g
QX#Q
�������㎆e���7W���[/E�Vg�PM���=X�Gv��<�����aҤR��q���a��h�XLI����UI�!�� ]������[��	�9Q�A"�ҵڠ#d�+�[��v,ӣZKt��d��qf7�va��fABzQ��_�ҕk��Mo�{��aDϿQ?fw��g� ��E� �a�<�R82XlxVHYEB    da59    2e30����~�?��L�9�9��Ґ��jb@I����|2MU<i�r(�gK�-�� �<v�W���F������,���`[h��	Pi����ܧ�ɏu��^p��>`W0|8���5l�����B���f��cAT������XC��K��;e�-v�z�hƲ#3����r+�����Ҁo=aT�/�36�;�+MmtE�U��Щ��hw��\����]BO�+ o��XDN�+kw�K��?}mդ7|՟GE��:��e�:ɤ�f���Yؓ�Pf�ҏ4�%��E���<���ݽH�ي��:��˚"7��4l����۾[I��	L�n�٣|)}&���S��(����j�L$�|X����n�?H�EvNL��ْ��C/�kj價ü1������t���^���6�<��[a7.)�f�3���5�������zD���&.;]���'p�z
�#�]#��:7υ,�Vp7*���!���~z�H�.(�m܁w�~��O_0�c�/dP���az$.�x]mZ�ۥְ֓>]�F49U|�@ː
��Q
Ji�a�E0�f��K`� ��:���@���mJ%���� ׈ݫ2�s���3_��s2�ic%$;3�v�F��vsɾ·!W=���#S�̅���`�9��IJ��ꮩk��=F��ưa�  ��N"	H���\�}��ج!�x�w�0�^��RE�*а��Y�ƹA'_
���SF�޻��Et��ƛ�(1:99ux$&`�$�+��1�x)�Í�������uQ����1hr��
H5���č�TI�j1*��1�뽉�./̹d��h�;����D�\�<��)ec~Q1�@�t�&�����7�\�O��f��x����@K�KT+�z�/������#�!�z��ܸxf�Yb��'�)3�]X�r�#��C%�*��y& �����v�|��2�/o~��@� nIJu�䊙���a߽�	�=�9��e��8�0���ld��r�'q5ޟ~��%��bN����@[�U��2��'�}
?2��B�q�biA�Fy�)�N[�pb�n B5q�cR��KSQЬ��q)���b3�����~�櫊�{|�����;g����P&IP��G�v?�@��A:�s�jBt�� DNˁ�	>���~ac3���~��骸E(����_4mҖ��t#h�����߂��]�3��������bDAyW�e%	V:d���	�䠬�H$��cK���`K]y5�&Y��Kkk/�i���cOz�ӑW��R��#N�$�AS���⛛�]�RE��|�ޮ�N�sd�O����MC㈁UE�2������E��Yqv+l�EѤ�װX~d4m)�7�wBhd���#�p��,��Gť��e��E�H����l�=�k�<�~�ATE�����8��b�]�&�'\��EF�DP�v�iP �{�-3v����~stla��<�~��P1OD<J�]ׁo2�����K]��Q�0�����_�K�6�դ��g�JR�� \�Q���F��>c�s�h�`а����R
қ)[�J.��xm��F��c��i5��Scš�OQq�Ԇ��ӇD��d�e	g�[r��:	���UvW��U��KQ��f�%��L��8��Xԡ؄�
�x��0���?){���y])�2�rs�v@:��	�7������u�x?`�'K�F.o�\
��츿�^��?����ϟ٘Qr*���IaB�S��6c/z��*g9������Jtq[��q�Ì�N�������!� ��z��B�� v7��Y]���Y����>sྭO��.�����<��ϼ�Y�o�nNd��G@�c ���� �pT�˦�j��<���*�|�QùY�&U@k{����J� T�<�r��b�ʜ��'`����kO8��܈�B)��eH��Fɼ+:B3����n*p4��>S�k��j G�|x��,����<����&pڣ�ΞW~��9X�w�p.��!B�
��U"'%M��;�wݷJ\q9��%�b~�?�E�$\�Ge����@�a�fwN�%�I��;FJ@C)�uY�ܓ����7?�1k�0�b)I;���ڇ_�LmoV�E>3Lr.W�J�L�罣����5�_du�OpٵK��Sh���U����"P�\4�;���p��d(d{D|��)�_܎�����mõsM�W=Et�rZx���o����"Л
s(�����?�ۅ~��G_d�f��G<�hL�7�^<��+����h��� � gk��A�̃%���&���͞�)�	�)q�3Sc]�(����/r��<�<���ǰJ��H��0C�" ��YO�� 4��+���D���n�k��m��5�P��m��rU�9ً��y��3<yL�g\�}r8-1�9���ٛ_�wa�&���"�問ph�m���N�˓=D�A��o49~Z^w62	����Ik�sӑ	~]�<��j�woϯ�m�W�:#�yR��%��~
�]-0���Z�FM������K@0t��١����e�K9p�⯠�D��ȲֳfxF�%�8��i*3��- }��U3�4����؏"���4�ށ�����O?�}�� 
�O��p����˰[�ۢ!&d)&�HG�~?��D�T���y�:�{EO�qHo�?���H�n��k�0�
��{PX�<���˨C�7�OC�z3�6\�vX\8����:�n�Et36E=���rѐq�l�c��e� f~�"~dV��KL�W4�s@�8��J=�	~y@��wh��������?���\��TE+�S���3�@��h߫�4( �"xt��E�M�*7{�u|\�GW�
31�I� q�V�}��Up�]�O¸YKQ+���wneA��b�9������MiG�Z�#
���"�]�H�,���`ƌ�����Z�n�fE}~Pv��Ck/��!�hxT|f�Ļ�m��BU�ڬY���Ԛ�_�/���a�qp�	�տ��U*#�D�0m�}�h�����Q(���3�{�I�p��΃��,!��y����4G��d�ۘEӤ�s9��k�5m�|R�/�g9�Ys"fJ�0Xe�=;�^#��߲���I��*[`�gOޛ6�D����� ��c�_��i܁a��1�N�taj6��"A��(-�3}P�;8����yV�bN'  ���L���5�l�5C��4?��;�,A���-���s�v!���Sp���8	4��/�Y�ܪ�H�ʪ6Ұf<8�0x�w*�7Z]���l.������sͼY��:Ũ���[��WF�8^Zt<Aj�pOכg���>O���%�,v���-�I˓h�]�fDeoK�Mb�n!U���~�3����y������pd��03�cE
������K�su$�T�F�\���tp�L�ϔ��`y����z �"(�wk��C���Cc�ȀX#K��!_ӥL�:��Cw���I���<!up<�W����e$3��l��U��7�~���0@׼�Dz��-u|Ov-0����#���1S��Tk�m��cDB_���'xM`�-�m�n=���1��9��(5�}y�3;L9N���Z���E���j���gy���i$ɳ�ʍ����{l6��jFM�{%��� ��r�ɽ����v�͝���H*���Y����+^�"��8�d-�*�A�= ��N��cU�P�<�0Q�5w�n�o���^�p���}���ˀ|6�-�{n�qI?�o��e�z�j@5T�#Ư-#���p^���q)��L�ک��Y�4[�y��'P��$��$5�4���|Lp[Qգ�-{����I����@�0eKֻ=�),J��؆�v!�s?���V��LDHR��sc�ᄊ�D�<P�&UQ�/1����6��4�jaхX���nJ�[��R��W����M�uW2%qd��Qz���'��	|`��KV��c�m�Z�9ob�Ĥe+������b��|�HOv+�ܥi0�h�/�R(>ݏ|��$��:y�:㎫��h���-��Z7�*�	�m��]�C����x͌?o/ T�J%�3锑a׊j�ф/yuF=�t)X�'�y�G_T�\3�sӿ�@�j
�j;��^�m��(\q.��=������̠3����lXX�{��}�tD#�Ĉ��{Y��9=��l:x?u��Z1���59~ס����������]:�~��Rf��ϸ��u�ڽ8����>@+��z�_����]�{r�؋�ӳ��+K^[�}�����@����<�n a��eh��F���Ĺ�Pn� �-�*f������a�$Og��v#���է�����Y�gl���[#�o��b��9�c%T��T��X���(^ u|6���q�����I��jKHo��1L߬d��}~�x��T��1���0��^�q�����Nc��pݻ�b	�?ƕ훊��eL�4���Z?���R��JG�+����y+I���nH��2C����T�9�~e�f�L������G�Q�'��W����������#C��l����˹K�XaГT�j~&�� �I�S�;N�w��Q|��� �5�Z�������U��:�e�c���1�t �4L�H�}�R����i&��XP��hh�������4�����L�m�#e�a��ޟ>��%���E�t�gwܿw|3m�&�D�@�ؔ�� 0��Q��E�O:�`y��GK]={}�'�r�pT%g�"���]�0��P)�ˊmi�G�]��;��1�Mg�����1�DŻ'�7�j����~�
`��>(E\�����3Ʊ0�N�ެ�tk�{���I		��!� ��tA�
#�Sg%��:�n��P%����IY㇜�d����$�0�٨>N�i��2}>� �����U컦�>vGó���a�}���� ��
u��誄���k�R�n3�_�%���v�[2�r*�K�	���3՘ ������	��+ܶ�/�x	��6��8xf�1a��E��M����{ D�7&`&5'�����Wx3����,8��X��n�TV�ʊ��{5e�WIQ�r��(x��HM�JE�iB�t5�%�#��Aϊ&��:��~����2����ڻw]�!ʈ�]�_rZ<~�G6���	PB�'���šM�����I(]l4�!���v~/3c1q\}�z����=�`�	x���]�<@M�~�����R(�P�NM����N,�HLИJ_`���SF)��c�
��ք���k��M'��!��r��.�S�>��$}��_ob���g�%��M�lH�5):Y��H������ݥc.c�\�'�.�7���Vhm3�\/��ʐ1!]���>]7�8���mW�qzC(�!�!�@�Y��� n+v��N,�iWد��mB���k��!�w���Y?��0�zĳQ��]'i2d}��wҙ	�'�q���+��6������f����t'��+�R�Q]�Μ��B�Q���9ô�y�h��C$�%䎵H�t��U#1�N�ٲ��{֏��y��'{=�O��>��"RG�L�T��� >"?S����Hb[s}����~a����\�/���=_.�lf���-�-����N0��G�}:s;"٥��x>

��n�O�<�^� )u����͵t��oH�0]��o��2i�F�0��%�EA����OS%$Rl���l���G�M@���nY;lo�R�h�xZ ���\�x�Z�e䳒'�k�_�vCc|;�,��?Q��qO�EJ	(�1�çz;�*�e����N���������
�w���_n�}�� %���DK]�d�"��Աy8�6�|H*0��u}��%�@��_��Ae�Y�׆]��O*�-�x�.2���2�;Q/wQ�Q�
1Z���5/ _��;�������Q�Q[���?"]�T�D82����l��`^�2ߑ�b�w}qh"~�D��Wp���*�6��>:L����H=b�@u�c����<��-ȟ0��OH����h�����v�u�b��j����	��I�` �$ۊ�lR��Bu7s���k��=��}�jx��a�f�/S���K��TG�E@��u�9Z�;����^���h7�L9qANC@�N�W���5�)+�I
���D(������
g&��qު��Y�7L�����me3��w�_wE�5�"> [N�SI꯷�J7�������m�݈�o���,+F��[`J���@�!��/{�%�%�[��.�wx~p}�[D�� h�_�$���Gݴ+�8�ޢ,�LOowh�1�F��6�!�ovŷ<o��"n����ܒ�i��Q�˨�"��G!�ZR֊��4�^i�9ƽ;��+2��1���.�sՄ/���!z=�}������^���h��? �t��q�b+Q��<����\��a�ɝ��[��x:{�3�DC�L�{E@J7z��@UH��+�7Ɩ�f�$�\(�ذv,o��W��0���A�څ���W�B�8}���#m���Af�9I٣c$�?�w�
�vy�|�T<�b9�!M6�yU�D���FPѿ?Ц8i�%�P�Lui�9N��`��iG��V䧭�tH��=w��t��w�u}�������W3u���|α�Q�_��ob=��u6��z��@��ɔ2�3W�yi���.��Z G�TZ�9��f~- �X�D����DȆv���	g{�iR��7S��-���*���Cz�c�ΐ���N�c���������u�����x͞�#CH�:8���Le���,~w8�j�����_�NU�;����z@ԯ��P��*�#�Y���rN/��-�}�ܱ�ݴ�G��`:�%h|��}���^��a�=�d(I������:����X���e1��&|P
����a�9\�JX�&�*�������D�#�;|t�L��G�X�������V�ȋ�eH��yf;�:�z�/xFl^�_}�Ә��g�&��B���ԓ��-(�;sv��4m��0�ȧ��T�M�NYGc'���2�7bW �Wzp�買��(��v��
L��'�uq���;�oW��,<���p/1+�Χ��>_vƏꋩӆ���W��:��J���J��~+�[��>�7Rr����fֆ%��OP/���\q�H��_J�����27�5��	�1��!o[��y'��Z��qN?���g��Z�q�w�R;x���?��D�=5N{�=14iœi_2Q��1���k� �n��Oa[�6����UBN6�8u�����+C`�3;���$��
�0���`�+[���k�u}G���l� �$X���	��߇���
P��aD�@��ن���
ON�,z�'&��(����IP/7ЦE
)q�k�O"�ĝGM��[zMtY�28��n:��svI����Ͱ�ƈ�ī��f�y�N/J�����ئ��~i4*��A~R����[j�4+D��R�J�2|}K,�$Ӟ&/5*�!����`�Lh��O�J�.'7d�wƭ�Z+�ɱ�^6�DZ����uC�w�.��#>.��5u���<�z���H 8�+��j> ߗ�g�l�YH�������U&:����Hy4���'���"M�/6V���v͸� ���0| ���VR�~<t˿���[�H�t$ӣ����!��z�[�)b��8�tl_ʭ2������5i�R��s�����37{&~"��3y�G�Wg�o�kݪVO;��Ǭ��O�v]7q��+�
k�M�.;«:[��U�߀>�:$pLl��s�ڽ���8��k$?��(~���Zo	��Z�c<��=Z��L".2�V�.�f\B�?�Y��1�#x'�!�}3�J���Z�D*�v�Tz)��T�f���lU��������b����B7Y�h#Цu;���PX�Ox�G�5�P�O�t%p)�t#���ƒ^������������{����>ؔ����	����#�a�0WMb�%�D�t������u<�{���-r�%�x��2
U�u�V�D�0�K�����)Ge� ѝ\��7T�}��v���v��Sk�r�gHK�c&��Ilj�'�#��[�_곥�ٔDC�by ��1�o��C'-����#�:Bh�/���8�L��Ĥ�%E�U�c��J9�¼pHW#-�WK�ո�:�kɆ�޴�/P���H�xk5=O0�[�������Y�A��}�l�#�sf�L�Q�A�8l�F�F@t5%T&%�;߱�s�-�fe��Vz����<��Df>\�I�m���I���{�SXT&"�χ����<�;�%�σ'N��O�����J
��=y��� E�8�2�EVr�\��
ʼ�F�<�A���Q��¾�K��խ���_f28��gS+j;S�@MM���V� 1��<n��U�s�^���$_L��=������d��3Rx������\���=�G���^����U|�U���fm���2��2�q)�!{-+	dL�GK���pyx)J4X+5x����UAZa�H�Y�BoQ�YS���W����g,#*�Y�l����e��#�Q��� ����9����^���\�����,yE~���=Z�O��;�
�� Ƞ��,qP��}�|�3�)���	Ǆ�W3��N�dcѕ�j�Iy������R<�*8-�+�h�6��?�#�s4p�U�
��㉔P��0�4��R��$	���{A����Nۉ D]���8d\� I���EZ������_�_�ɞ��%벜3;�R���RJ"����i~��<�x,"ƾ�����z�������l�<�R칮֒���m���М��@�g�Kz��F��F8�S\��޸�r��A�)4\�O�v��v�LqINajؤ '���7ar�B����~�D��A���j/c��n�'��:��Gɍ!T������&G*7Ru��j�V:F����Ӥ	�_I���s�]����@�%y�޵�X�;�1 MH��\7���f0�����(����Xp��Swz�ʉU;ɱ��qdZ����Y/��bjzOR�b'Áʚ| ������h��B-��M8q>(g	����*9�B�3���v�J��ߑPڔ!���Cn*��0ϭwot�'Q6�i4C`��M�GC��Y�m������BX:���l�
6�8���}Q���C��q�E����ȱ����6�ܯq
&;Du��Q��D��<hq��")��r�VG�Pv�'Z�a`I$ܔ�˷���1p�㓢�$iZ6{_z�wb�\��
�{sJ"{
� �0��@�ݬ����a�}��ذ��̮�����+�2�\;ޞ�Џ�<t�|��f?�<�Xn����]'���K���Yej{��ձZ�B;��-�8�J.��!0Ď�j�oaY"��"�I���,|.��AQ^/������1Wt��) �E������9Κ�\�U�e��CZKi��#�!�;?���J祠[E)j�a>�u
z�z[C.�P��=�b����b�=�X,��+;�o�LP_!�d%+�#�l�*������.���Ԫ⻉���{)�.9��L ԫ��}6��{2�����g��F\u1��'�B_��;hy̎�#����j����J��E��ѓH���D�j�ҝ g#%67m=��s�fy�}�_m�ߺ@�OZU�a�� R�E�M����f�n�p�4��\�V
�drTJ�d1�K�2P"P+q�����Nu0gJ+y��K�s��	�����#\�����;��S���"��=b��δ�ś��//o�4�=l��Yeh"9윋~Oq����0b,�i3~L���)�Y)� �{%5*'DEJ��T�b�F�&&Z�@H�����g�鑮;xC��㩈6 $�n~/��X�=}����km72���E�P�	��D�B�R�A�a�C�'4��r��?7�$	b�?������Gƥ�D�Sf�pz�+X�io�`��4)��f�����kyd� }��\�u�����B��)|�1lb�}
�R�[��E|���B�����
���JH�y=(�����L���$�M
�!UL��/�����4m�"r�{���?�#|�b(�"B�	�CA)�^K��y�3����*3�A��z[{�K/m�����2��@5+0�N�*�A�D�5���5����c ��K����3~��.��D�v�Wu�L����gX-`�ϳ������r��_;EWA�<NK��㸪�O��1�W[�۰[}8���݄�]�Sr��
�&�f�|�I�tݸ��0z���@��=m�`�#	���ц۱�v�P�[>�kM�剋{ A ,Q83����N.��C��ט)@i#���m�0�}������X/��1B��8�8}��Nh�������Y�1�lH*N�Z�|]6/�њJ
�pz�¼>tJ�C��䊒��������Fda��<��IA����"dT��'���Ά<�V��6�l��UҀ�o��p�V6b|_#�x� 6���v��守�(��R����"B�LN���&I�z��m~j5`cb���:�62
f�
I� �H�e�U��$�Y����⚷����$a]��p�1"�^�N��N9l��Ւ^p ��*pD��Gc�ަvb����-�1c���� 4���� �]���<��i�e�-P���|!~�:�'4��G��$Zu�犳�5��l�� �%��Cg<���:��>v!Hv�=Q(��ǡ�V�Q�3t�P
O2�r���?��cZ���NP^xg���b!����ĀFbI7�۳���@ג�Fŝ����FL����޸�DYf�IA<S��.\nJ�6+�����7+e��CW�>W)��@u]j�6z1�����tI���x�ࣔ����~l���QZ��}�G�!���Ղp{x�ө�5�1"�B�ɀ9F*�2�O��*�մm��F:�B��R��/�����!!���0j`�ջþ�Q".Ԩ���t��ő�U��=�_�u�S��a��,���d�� �R9�E����I5U��q�\�PoD��Rݻ|Js�0�n#t�r�>�V�Y���G�X>&�}P-j+1�B�U���|���AV	���;�3ҟ}���d�����>��h:p�Yq=4_����?�zb���Ѽ/�,��2R-#����Lr��X�_k�R�򨍶��� ��3��.ݴM����|\�ڟל�%}=7���L��d��wP�'��g��:��w}��X���xD�I�kܰyÔ�𠈬�P�cK�7�Ҫ����_�����3����s��J�H�|o�(��K4����2���y�D:���G�=��F��{�(��D��g��h8;y"�?�~�����«�ܐ��r� �TP�L����V+|Sa��ʵ�|�.|����ɷ��ff��ٓ���v�	�k`�*�J��B�>^�7��݄�6y�Qi�
�(v�%����u��1��#�l����Ѽ_&��F�ET���5x�$��w��;�i�f{��d�䘞ݑ}�|	�Oh�H�� rj�G��ō��|lk�,k1�%�I�r��єdXAYY�Y^<>�^��C��t����6�R6�S��:\	k�\6[zed-j}�#�e