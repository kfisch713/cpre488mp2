XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r���0���)3�:8#O�I2�@B�Ϧ��l���T�'[A��{�OC���D���%�D�����JS�h3P9)���h�����-�&4��ϭ�k�j� ��m��j��M��tQ?3�L>�=�O�.�~Fr�F��[���o�:\+�>�k�%��hBJ��(�&IVDZ����8U=�Kv���M��i�MQ���u�8��Jb���
����6U&��k$;]������,�"O���Hv�~v�/�l�����ZO0c�?=�[�a{��2���Ӌ0vG�"`Ϟ�����zJ
�.	�k��#��-'��ސz���o�?��',0��`��)sӺaB<�!�>����)6�p5�?�k�.w�q/Y��J��A������g;��w������xF/��ih#g0�S����Q�]g1���3�W(OS���� �[��E^8�<ӼB�?��D��b��v����\=F|�#Z\Q�9+�9츀n�w �\��7���ɂ��3�/�a7��ߏŷ��9�I��H\Ӟ״A��LL�GU�ٻ����?��uڬ�P�����S3Y�n�[o�A�� �'��nX3T�S��@�߫��ڄ&�R��h��m�7__YQV������Ϸ��S��Sj���n*�m��,-��qIߔ�Ԓm�~�RI4iə^��] 8j����,�����J�%$c|�[/�Y	y���7���&M��ŀՑ[��e��f�Uv`��j��!�4(_��N�:�XlxVHYEB    3b09     f80��?( �Չ]o�l�&a�<v5��#qu������3��Q���ہ�1���jk��j}� p�E7t�`	�q�f{�k���i�!H����F(��@Jp����Z̈́�F81h�']0@��)/��H���`g�1�֔�u�K��`�Nb�=̫i4�� 6�*����D��E
��8���Z	����-�<���[�1)�!z@-��`�@�;%tOu�ږMC�v���)��!|}��E�HT:
jFv��.����7���yH�R�<�$W��u&�²m:���hS%�)�9_F�ųB!�lf?�d��O*�^X�nߴ���$���%ߪu�L�Ͽ�d�ͪ��i7¡���d������Eǋ( �vڑ*��.�5F'��@Sܰ�� �?މ�gb��_?��p�^Tu����sf@-i
a�Y�����x����u�`��\�i��^:���o����Ů�33�@��\ENP$羿��n�}�+3��Σ�98����:�\٨ÛbwvN5��&�LVꎉ�Fb�츈�� �Ԫ���#Ɵ댟I���
;��z��"?���7�L �
uѱ&~�ˠ��G
P�Y�G�{@��&�(��TG�9�Ǽg��Ϥ�r\�'��8�T����?:Ի_̍�g�$��L��*��f~�͒ا�I~�=�,}�c�F�dC��w�B��N0ad�`�^�K��.�J�'��)l����:t)��^�uu/[�]&Ɵ�0�RXK�!���,�a�j�"�d�ܟ�y6Z��[�7(
lː��	S<���;Nɍ^q#_{J>��q��\Cn����p,�9�ds��t3YR���W��]�F�R��[h��n6�J�)|,�;W3OV�҇��#���,*'$>��6��dw�*Ӫ���;!-�ԣG:��qٲ�0�����z��B/^^'W�蹗���0�9�N� J	���1�ƅ��[:~������<5E?���h����N(w_8S5d��D�d�Ӧ���>��.T���`�?Hj�@x/'�2P����|�;��B=�1w��U��ص�ʓ��/�D��:n�e��U��~E�g�`�u^�Jw���|����ȥ�RCr��fH�2������au}C��XC�	�!�+����Q3�d���	Lk��v>��A��:G�m<I�(�U�gcuڣ��y���/��O�1���t��X��Ȋ]&*U���ܯݺ%x��G��l��\|4�o��±_Ӽ��Z�v�_&
^Z�V�^���䑊����\w��߱OSuG��zo��|�κ�=U4~���
Uu�����[#��$�3��8B,�'�I�aۿ�,����n7������W���*Pq����V�����~('^p:WZ��5!d�=%�� <:*�����x�f<Y'��+WJ�tdGݴ2[/b%���	F؇���g�~ik{�&~\^��~� o�9UX��\���5�½��`Eb좺�� �����V�����Ds��:����tåenG�Y�XX��[�u1Tn����5���
�{���567 w�$�K,�+��ʿ0i(��0i��>�f�`ڝ�ϻ��!��*6)�x`5ri�2��7&ÄV^bKh3��?��w3w6���B�f��'4������Y��o�nD~v?n��DM+�I�ϯ�3�.iF���k��]�*�`�0�ݎ���Z���LR�����e�`��~�B���FԔSW���,��o�K�_8�������G~�@T���K߇���ӥ�C�//Ng��i�%����#�&�^>�2 +r����ĺ˽��t*�@	/ŰΔ����J|ٺu*L��~~���K)�[#�9�E��̏�{�w����M=N��*}%�J٬/����J`ݬ�8@QG%�W�(�ΟM�v�#�PCV�| z�i�.���@HM�}��z���qX+�TuB~�ѡ��U,��Hd@O�KF�?�X��!���%K�N3�I� ��迧_܇t��2�F�I�]��*������Z����hd�K�>U�55���&�����v]W�߸��Km9Z�cz�k�O�i���it��8r`�E04�?_��d �n��y1���_M����w��A�<ˉ�7����f2���C��c�_��O-`1D ��D�պ#J�4ۓ��)�6{�w��y]PUt�Dsw�L	a2��^  ��z�Y]A
|mIbM;�4.�������`��B�x)J����V�E�7��4�O`CEJ��0���с��;��]���*�`�?(o���MuH�ŏ��k%�A������|�3N�wj,��M�7GY��y-(Λ��RV�6�e�fLؽ��d��xϭیD���}��g._����N����d�^�����UP��h�lG�W���2n5j��3q��}|@4cׂ��ᕊ4�@{��v������K��A�W��__�W!����e^��d�L�N��ϯ+�y���A+�\�j��F����(X	����Դ�[��<�������I��c?����������l�7���0-�����~�+��1@�ZV$E��6�s>7s��:�u#�0��ʱ�zy�|�f�i�{i��e�5
FF�i�TmQg�M��uqʺF�b<�@�$��u�2����ߢ�K�.&+���˧����'�^�jVS�L�Z��Cm���Z��ٝ����N|���'T����V�D�����kE���1�rtHB�诟�	���3 ��a��0�v��<���K����F�;H�q"BnTۊI�{n��k+��Dc�Z]�EG�'2��"�DC9�_�s
D;�������2f^�����`�Vm<�m[���^�x(>��%�=���l3���"��^����׈����-G�H>�1�ׅ֟�+C����k�|9�x9��T�Q���N�ŏ��6��F~�CA���w�1�3X{�lӞd�5���k������.��~v��]:�5o�|��QN��g�+�n�&T�[F"^��f���(ݖ"LZm�Et�ƺ��L+Q�W��:)D�~���1W+����	M��?��\�%U�g�k0N���t���b��_�9��?�9E`2��P6�d.�~�fl��b���\`�?tR�R�1�,�x=����Tz����Y&̀�u�fS�E��AU�g߬���V^���}���g#��U��t�����:�\��Fw����lo�3as������V���M���V��kT�E(J����4齶;r�#����rpB�L�*��p�5?dg����LRږxn�%������Ai���9�z��� 킆�J-s:i[H%.�U�~�J��P+�H������e��1*�VYa��]��%ð��V�.{����)�28=�(М��ӷBVS����̧*7�Mp�,©+���!��}��kj3f.\�Nx�ꂰ�!��E�q�n�1���'PзCn��=�s( �f��/,��"�;��2��O��?�y��+bO�0�{�@bn��"��F��
�����i�sg'���J�^Y~e!T�=�^��@���ݝ(�*��='�ˍ!�u_�SXX@�컿�p<���|��s4�z��wP��&� 6^�5?Q�*�Sr�aR�!\p�����l�c;�(M��J]j���*g�1��g���ǣne<&q��v��~ǌ������p�ҼKp�I�F��Y����\�P��1Z��������}<��Q����M1=�s�M�]�S�puۛf�>�	'c{��Q�z�u42��%����_7Eʁ-Lp"�m6��ݟ� KZee�Z�3�X�,	�(BqkC�}����h0����3�({0�ObW��8i���BvL�w)�*��WG뙧%Ǐ�e=���͹=