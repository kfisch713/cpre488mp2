XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�P��J�0!����Ej�a���!ݵg׬^�M1\j�9��������c�/lǬ��~��A�+�1��J���ANIm�O	k�ޢ��Y�WP�.�rҽ
AbCў5VF���⎫��2޻�����J�����6I�̯���B�Y����ڕh��I,jd�k��٬�-�,,�YZ'�;�6���� ����yC%�]}�������\�yd��ˆ+җdm��H�E��Kb�ۅ���U<��T�g�W5�Ӹ����9�V����&�`?i�L�]jZGM?�o�X"B��d�	�c�q�{I�1(������<6���?$�����b\S�]�_��n��2�Qa>��St��7P�ȡ>KYd� ~��\�2�oր ô���^6�G-#��A������]�V̕��ѱlhj�����&)k�#��^��vкL�w� J��T ���E���o3�Aۤ�hg��X��_z:��x�j�D�X�Y2/�Fp�4�j�]���A����O`�b�w����.�6mt���T6�T���[���{��ӏs.j&q0��m~�a���*��L2���_X�]J^��54=3��x��� ���_}�D��+{jch�ê0 ���ke��y�oi�W�*D�iM#�$���^�����dY��L{���r@+�e�{��Vس�7�Ӡ��c�����w�a;wr>zOIY�6�h[d�7���Z��ξ�_���]��q�ډ���S10r����8mXlxVHYEB    5fea    1830D߸X�+D.$����c�������@�ӳ����e���n%��n�!�,[�(
7��Bϝ��q��ma�g�������̎Dw��y&;C�����D��m^��v*�B��$Fن���T�v|^R��?���ZJ�XؐGJ�p�������zID�,o�dp�V^S Ίn�it�W>��4�&W��Ǟ�s��'ZG��ݿj>+����o����?t/����:�#��zxф��E;��[̟n�Ad���h�h3����i=J�Jk8���),]������N��Pg��[:8����	#IÓ���ܸ���;���11s=b!�>�ȃ�A�{���+�]�wY��cW�A`�[c;�\�"R�O�9���G[0+`&��#�%���|����N��o�������г,mʲS��ޒx�!Y�λQD� i�ƍ�k�+:������M��RCYk�ZYO*"�A���b����\���M�I�Mg����C['��/����� V�6P7�_�e�y.f\+�����4:L���EDɬ��d�lt�h�3�3��HN�ȷ��v�0�6	j��{���&�������Â�]q#QӾ?.h�Ԋ�-Y(�N�����
I`9��}$�=�6m�.�ޫTft
��H�&�q�N�&�yabXˑQ����;�vؙ�K	���GG��4Z(M�O5`�M���	&��J�VD��;�q�r؎�[�[
���#�U&	���yas�u�7Au&7!Z���Y�d��$$A���a�A��J]b�u������Mk���Kt�%L�@ό����T�9sw*H���Wel��7�#<���^�
P�b��<�ı�gб��{8�����\��k�`hT�/s�V�}E�Y3�ތ�d^����t����.d���0$�y��8�h�M�/������#����sD��+�>V�^�������pM�{-�$�
4���V�M�5��籪a���"7Ǖ_;DzGGDZa�h�r�
�a���������Y���6��6 �0@���
��B�/�q�#��
�ct��k���l�O�KH���z2����2Ķ�Aˁ˫'_��z�	���x�wx�� G�
�iI�NgB9���P�n�w����=WݕZ�45�xo�[ɍ��G(�{���}V!�K��-���	# 9�d;	���`�
��H�Jd�;O�Fx,�Ld~!�/�5�31�㎈�[��jz�k�+�U��n0{QBK�B�=�����Ƈx)^�T�J���/ʿ^�J��>�\��|��C��$uE`�����~�v�[��Kf ���v��w�
�7��42'G������e�?y�ۈM�z�nID�)��-���W�;ͻ��-��e����.|1J������ɠ(bg��Q�\�5�A���遁�B T����LeC+&����1�z�O`P���x����V:%�mXe����:z�����M`�$�sH�)M��i�
���.����8hާ�_�j�ʪ(茠�(#$d:��'�펃
~�=�? V�U8��h�F�7X>�Q��X��]Kց_ݢ�	7��f�:�|����+�\�7��eNxu��W8
�a(����3>������?��^���уq��mEb����tNEsy����zK˔�l���X� t.!�|)����SR�� ���r6���#m2�2YHQn�t��rW�+izo=��z qv�`���
z&k��Ƀ5,#5��!����ci̓p9���K�
��+P��XR�-e��g����{Q䴘�f|H��T�q�_�lp��ڲ6l�a����_S�ŗ���V��ѣ�}[���S��v��Ё����F4O��Βw�m�X1���-�����R�;w
QR�n5�!�{/��9\^.������k�G��6�`q��`�c,��B�d)�gH�j��,���i�-��)���������@�%s)�b��B�4L���Qm�y,�O6~{��4��p�ӨƀYp��0������n^�CC�ޛ���{�ߋ���ΓF�@d����&���$��	g&�����l	�Q�/��e�ݽZA��߲�k��+��O���BA��B�������B=�`��*/���_�`�-N��a�I�BU�i 5��ֻ��粴{�x\V͜��ܜ�2[$����8u� �z�}�	ǘ�fC��B�I��r��Ȣn�T�˳���%!k�����j���V%������_��A��Cu����yO�T6l�����;:R����K�9d�zb?!?B���G���p;Vu�X��l�Xe�	x)��y4���U��b�̺"<�h��z�B���b��c=Z#�*��	´�*|w.ݬ��E���z���O�\a�6ޫٛ��
PV��Er�~,H�x�v�9�n�F��!H!�W�l��RE칾�!��+���?���g�jɧH��4����L���r2�|�;�uHa��	$/�j�@��nQ֞�@p���J�����T-�e�
"��Z�r5�q�&�6������H>Aہ�:�0xZHɌqt�|d���UҬ�k�E�́+��5v� Y�f�MFl�-��ӧ�k!�.�zQ�at�Bd�Զ�h�_>A�%}bs8٢�SM�2�hۮ����k�L�.G����؞Ih3(Z��8���Ma�U��I��ѐ�C�������_K��<c<���:��B�v�P�c�*C��US�a�J�]PB�҇�����r�:6��a�[��ȹ�����4������G܈�� ;~LpW(�\F��DS9A��D�{����{��7���I4jv"q���_C#�;k<�v�,�����ف�����;�74`5%��}��$*�p��:!�.�+k�`�L`<�Pi�ޑ�w�id�Py=�������>�Oi��W;��kNr��-��C2�/�֓����M�
��P����"�F2�p6b9������E:�?� ���D�z�)����*�ׁ�,<g�f�~2|I��~�vP�n�2罎Ntg&���o�i)u3��@�i���K�f�!��-~��נ9���5`�$�>7��j���>'�ʚ�-P�#�]�>���#�l�9���t�;P�jB,�uﳒ��,K�Ja�$6q͕g�ŁEL;�����z �+�.@&J$`I�̌m����P��q��n5�'�V��SD!�l�,�oJMϔ!�j8�W�\ ;�)��]��nt���)��}tp�OY� ��`�g�r7�<"t�/٤F~��v������PDJ:_K~�c��T"����H_";����!����:�r�#Y J�2�`�`�rm�����+�^M�BPnUԹSC=��Z���v�z��E�g�M����$���c�Zt?Z��Ca�[��T��"
�A>B�;�x�i��1��5�K�m �q������<�4-|z��qn9	���#���/����1pJ>�����2.*�O������F�T�Cw�+S����Sf4o�@^!U�
��](,�QL���m�`����4ȂT���k=1�22��w��q��(�L�[��O�*���9��u}�q���0��MI��i��+�u�§�\)�kH�&l+X��.@T�\Wq�HO +g��+��9ũ�էV0���Mqp���r��Ă;j���.nRԪV� 6��0���v�K��߼�O��?����C,��d�F4߉u�2G�$���Ew_ر�/;��E����9Q�����6/�E�t���x����W|�Y���a1���}t �g��`��#���������mY{t�#G�c�)��7�r7�����Ohyh�NU��J� [8���,r�$�+���}1��=+#�YE�5Y���B�Ҡ�e �ܦ�f\$����x;��W�W4��rG~ވ{).aͧ�����M�;��{�ay҇��wgxy�2>��w���lN��ͧK
��ަj����vj��T�s�g��G�� ��Ֆ�^/�s��2oM���bT]�Mӽ�I�<htu8����XL4�F-��flU�5��\��:�U�ז��g9\�J�q$�l��V�|�F�l&/�d�d�{����4�BXqLi�6À�!I�W��?Kp/*�[��a�N%"J�J��Jv�d�a�FYp�i硍:�|�1�m��_E,���3GJ��;4��я�?��{3K���%��"o��\ב�j����7
Y +��;�v"�9��I�ة*ؔ�܇�jY+���A����7w��(L�>�^�d5`��u�Uz�ݓ	���{/n���)�M��0;	���]~��Ly����,R@�T���n�X�|��/���C�����V{f,L�
��'wl�%Qy���_��5�c�G��Z��G��\��J�D��ô��jh`K��~��ե7Ь�R����Hj]ʒB�i>3f2"#�m?����1�6�I�mVѩ��|�8g���j�7��Z����о�_��ԹO��2F�?��oХ��o�S���D��\��&m�&I
1���ψ;"�]���9��y���ڪ�V3o�*��HS]�7��q��SNKA�K�A�[���J�e�1��:��z���V�(^�ꜳ,nK�I9$n3RغR����f���A�,8b@�k47>���VE�`+��ETvK�_��
�N�RG�q�y/�4��]���X�t���Cri�)[�Z	�7�D��pp�ヲKz��:u��nq�N�^�`�R] ���з�@�d�:�ҡ�^���,|��k���S�'�y��LH*�0���DP��s�M�'�Y�z`�'"ǧ�"P�R�3�隟��۪T
� J�Q�4�a�f��T"�9����$�u=�An��o��߮���$]X:�6��6��y?�6� N�0Wj�lJa�?��ɫB�lzJ3��b�j]�vx����=�~+��
�)��t��O�(P�Uq-��~� ^RӉ"��3)��A�^�vi$��Ǖٽ��M�z鞟�U�=a�>:�M������$�s�G�oj �*�1�0������	�:� :*q��o���0�絘vUd�#����Ӿ��b�[?Dw���M�",D !ͽNߺ�:h,�9�[�Ѧq�(�y�J��Ok�PGSM��E�L��N_Nv���gJ�Z.�@q����2i�d8��J���6`]
��8��k�0H���Mެ������?�s:�1�⪽;��g��ܤHN�P�D��5xv�H$-U��Z�����K���(��S������	�k����m�tsI��e0�n�����B-��ؿ1=�Y�B�����n[ ����$qEZ�!s������7Y����_���Ǫ_��R����+�@�Św�~����W2�#���NL��&D���,�I�u���a$cjtߥ��7����z)�=�b�17�29���׷4l���{�������B済� ����[ϴ�%'���q�M30Ƈ��(�;��}u��������DS�U.o>;�rx����u\(�2��Gnd= b���?��@�t�P�R�pyЯ�]g}Pc/K�5�u/8f���`���1�ɮ/�R��LԎV��U�Jr���ۓ���\Xv8����3��I�0a���_��[��\.	C\���c����e4�S�H
r{� ��x�#7����\eP �T��,6�9�s�e�Q
�iIMn�-|ܼK���.�y���w��k6Pg,��ʵ`0�������+7~�����"�Ug�@��=��M����Q{�@9Bn]$���ca���T20���[�;צw:�wXQZ�0dvš��#
Zp#�~�q��U��k�m�'�9t��i��ѕ��B#�Y����6o��������EҠ�4=�s��m�L�࠯�j����B|aφ��3갵=
t`�6얪�P{R ׈��Ɓ����5�����i$ZK��y�9��Z��^�<>\�M�dF�ՂƄ�h�I���5�
��gꛪh�՝���r�A1���0�<z�9���`�K;s���}/�|L��� ���df(�������z���,�<��+ӓ�Y������ȉz��o�BeL�m!c��������