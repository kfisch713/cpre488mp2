XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'�Q��
ۚDZb5t��\�:���2�v��O�)��(8+ɓ�˝�oU���^1Ԏ��F1��-s�ܕFn��sY���^3&$U�o����Q��֥1AVM���P_����p���)�����N:\�T\`:��Vk78�Ӆ?��E��K�ܷ�Μ<7O���=�0�^������i��ec.D;Q`ln��@��9O�ҁ�_-|�����-����Y䡏��AQ�'9/+;�=AY_J��M���^*^�Ƕv��v�s��U�/��1}�G�C�~d@Ul��7ޖf�@��d��˦������5(�Q要����X�%���'M���@5�i��.Sc�������`�;�y5��8��/��-À�ٵ��W�(X�����xm�@XX&E&���/�w�6���=)��v�i(��@� ���\�@���o[�-&�J�2@�s|%N����ZG��A��~���B!�o����ѡl _Z��J�-̾w��e�S���y/���V:f�����U����;�%��Lrt\�iJ�t(笐����t���2	 e�-�:
q�p͋�
P��ЙI��$v���P/�_&/��A�{.�0���]�|8|'�$]�iYm^mz���oM�Ih�M�Y5�sy�O^G��Qxd��ZR�/�_�����~;���0(�M0FG�j���M�M��jzX"̓y�[�Y���,����m��gQC>�֓�u���#�_[Aj�9oifZ�I,��yXlxVHYEB    2b39     b10X� >B0�)�Vl��Ա�ͧ{�P�P�Rk��^�n ��ݒX�D�I��$;8�*�4�fY����$�W��/����X�do��Oư7�z+ׂ2w^����wB�"�w\"�<���%R�A�Ur�Rj-�H-�"y�[�e��o��f=���¼��ԗ�QWY�b��~�nHlۮ�wI��n�(�*ڟq�b�g�՘�}y�f���G��;�p1�M��f�s�!���z]�� b
l�X#s7źi��{w�]>��.�6�.zZ�J��k�҈�`*��>܍��f�G-U=������1.�{dK	[滇��r<���<\�k�����M6D>��W���z�q��Ý�����}��ʜ��x�}J^^=�G]݀�^���YK�	`pv/ ��dkz���O��^F��;!yK�����̰.{pS:���BC=�f-1��
��UB�FM�g����P��S��Ǻ��>;�扚���uR}U3�S��z�D��zJ� 1��g˴�כڒ�Ƨ8�C�mǚD{F������ػ�,�g�Qc�}�Q�l�B�:������~��Bx#!*�\���>*4�X��i�m����*T�&/:cq���E�T`M�w�	p&2�H(q,S���=�<x<�z�$~f	[�o^�h4��_��Z!��e�P��v���~s�Lc��&,�s߿�'�����S�%��!3�zű�͎����	 pj��#D��N�k,)W`��&�����ߵ����@9�Ս�*d�#٪O�rP���
ͽspW�15ۣ��1����Ή������I{��!c�r��񣼀E��|����z�'���tJ^��C^�Q[�Ȁ{���R�Ίg��eh�����(���R�-Ij)G�s��;z3�>�C��c���&�'n�-�8a��
�DA���V�u>�#�5D�HE�E�r���X�h�4����|^:�����&X�D�!��.��\�9 �X��S�cc��y�m6I���[x��r�t�-;�O�s=w���F�E����}5��1qkHJ�,U��8S��'����f���OM���t5���H;��h�Z�"�$�N\<�}�c�?�zt�9���=�=�R.�uq���Y�2�� ��|�?�|�b��?Q���5g���� �}����x�F-.c54��i��ډh2��9�F���G�#�y��<Xs�'�usS��!z�%�b$�k�]l��>r?iA*�yO��}�ͅ�<�Vf�/_��#wյ��P��A8�SN1�O�����e�ϖ?ᨨ:���!fǐ��nNl�`��xs��P�ʉRLl*8٠�{�׃�K��0>�UC��2r��6���u\��T�+:�ߠm|B��S�B����`�o��p�_�!��<%���W�S�ɩ/r�G�Ay�W��a͢S�t�Y8�oS���]��iH�Hz�!L��ө�ꭙ:�G���Bq��͟>����@�lC�L��X��	������B5����
���c�Wl�r�v!�.R�]^2ݤ�� �7���f|9d%����Q�l�ee��2��Aqmr݁@?�E�O5w�!��a˸�o���>��}fH�3��ٞ7���q����K���u���?Pʻ�2F7{��٧6rwi�R��oE�j?�q�"���SyTS=_'������=���k���1�^�ւ0r�̵F����'�Y�ʄ������qS����=�n9��g�t�#�0*`?����� �SH�D��TP�Y!~}�3t�O7QQxL^�����+�8�Ϟ�Z�Z�h���,:+7dNsZhi<�R/�q��<�R�|�ѣ����U2��ૢ֦㐆���4Ǜ��Ú�&��[�_�u��΢�>˗K�Mx�|E>eb����{r���M]=r+AP�gb���=�[���I��� ��P�A�}Cg0�G#g_��P^��j:~�����m_k��tEc����IAv:��`�朷��H�[���3ȥ7p�{��酸�~5�6���z�C0�hݷ�U����'B?B��-��z�������.�}S��Q�!;�L�-�Wz7fNN|L�����wK���?SdV����Eh,.�nX`���L����f�Lm3�n��z��;�z��t���e��1��(��z��f��u��8��$ ����])��Y��e��,&JU������r0�]#S���- 7�&��nz[�~��(Up�ðZo(pݮc�Kֺ=z��E�����"z��%+}Y�u��=�3O���Dy$A�*LJ��=^���oPڞ�R��9o�H��ﰋ�H5���^�6	O�`�)��*1{����@|��X׿���v>�E0�v8��gX/J�DͲ���M@Ügq'�\��2�I�J������/tc�f�w����@u4��*�������nL1��ܠ�������0�����oީ����7��ad���7�$�}՝M)��
Tc�`{��]+؞�M�"���t2�0Ņ���d�P�n�������>��PΓ�_�jXN�|�O�C�0j���^R����Y�6��ըS�E�f��Y��\���6z�O��w�$���@��>(���@����l>w���J�4�7�X�qR��I*�~�QU��qh�%e@ �G��QCMz��tta.���i@C��o��l�n���R6��X@c���Z,ng��y�H�,W�;]������� ��I�m�.�Vx�v�!�C���#t��3�qp��
kj��ZD5�M���ֿ��	�.0�>zyA��J�X��y�B�3��Zpq?(H�T��i(