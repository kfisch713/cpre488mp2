XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$���Y{H`\M����H���a���@nk��EW�v�o�^LRǴ�T U>m�6@�����:��@��� b��zbW"�s��w	�>�p��5���A��=χi��ل��/y:c�8W����}\s����Y�ů�e�D�N�"�&|�α�ܽDjc&%���YԴ�k�4���
S�P�J�GsCG|p-簙�c���<7�&��{ڿ�qh��3�R(GŢ�e����&m�vq�4���ݶzߏ{g�ї�M3���U<�y4���N��Zʛ\x��"�:�&c{���u�_��<�܇U҃1qrX�Gi�%`���r,Y=&:�]L�o�,��?*o�c�ez���?\���%�C �K�M�l��Oow�5���<Û*k�bv �]���f&�R��xR߅ڒ���5�C@��j�ƁAJ8��"<�@$v_t��n������J���:����������>�6X|�br���}��k�n�@Sب�=�+�iq��B[�zdkmLoEI��@��HձEtٴ�/$V���A�z���ٱ�@3߭9�6ݒ����^^�*���i����@��H��l��Hi{�um�fu�a3k��?���L@)BJ�c���LG�h�zj�*Wd�N�J�hS93)����R�tCʤE����wȚ!S�|.�)[7������W���ι>��5Jm>��;�"~�=�Ô-���\0��H|�Loh�t�������\'e�B�A��d��u|�ʵXlxVHYEB    39de    1170y�bQ��n<O��㢿�)i�b�l��Z���@�ĸ��xh���3��?]��s�dLb�%a��>�
q�l{,j��X���a-�l�-�p�C�{V��k+��5��$*cGu���Lh1�X{����q\�PH*���*�-s�u�t�������2�	���ٝ���c�]4�͑��q���"Y&{y�ZO�_|�랙=tHQ	|J�dq�g�IɿU�|�M�id�w�0�������gF E�4�����q3si/ڈ�k���P���T}Ǆ�i30Cle20��bI�����$I�2ӎ�L���L�M��l��]F��"�.nJ�%�ΞrQ'�ᩲ� 5���<��E�f�ִS@��ߟ]}�s�����A�*#�\�|^�N�Д�t�-�tO�Ft���.z��$!Q��²�G�eD)A�hg�j�����/:�����X�;k���p6`	,@?��.8�rXHP�P���	��kڝ�d��~��6��x�!�h�aGn$��n�	X[��,*��L�5O�� '
c��cxK��\�A�n�D;�����!K>mE�`�K$*����B ��ᕷ:y���b��^8z�,�z���,�EU�H�u닜�9�����DXK7o�	M�c�pUdd�P� ����јL���0_�	y�s�˛4��h���2+"��ý��rO�	��R'�z�M?�pA��L�y���_���]���u{���%�Nu�m���|eh��7�]į�H�y����}Cm8�V����8N�ޙv��������i�	��XNU���.XK�?ݑpqM��z�E�"���,���]�2���:F�tb�M/�T��	P4�sv�f�r
g�7�V�s�+��E���R�j�)�����
#�P2�P�8���\��g�؜����09X�o�Q'Ϣ�n��e[�7Kw���Cr�(�P�0�c@�
��$�����d��T�)����g�� �?��,�𻲍|	�oC �t�q�A�G$��v��/���:;(���~� �X4�F�U�>�댿���7i:��jir�R~Y
ҥ0<F�#q�R��X�4��'�INi��L�v ��UXʉ�H �NK�@�~uܔ�A^�����;V�����v�M� -��ұ�Ns��B��xJj�ՂS�U��qgz^R�O3�ka�=�HPՓj/¬K�4��^	;~��k�JH�v���F�p_Ԁ�b���;#�m�k�FV۪O?���`�[�:@�s�H�u���6SS����IXUW��O<�
���܄C�Rw���V#I� ��,bkd�H	�U�(k-����(`W=�V�.ž���'�TQ\����4Uf�Z_q)�gu�-�B� ~.L�ohȂ~�hԫ����p�6b�ɕ�'�:��LOl�v/��{N�_u�oX��:�ld���!������	��Ħ]U��/�V26�_,<� v4�6�^ϧ�`�Aw�Dxe�O׾����p�KYA�Z&�����m�wZ��]TN�l;�Xp��2��}5<E���zxB�v�T�U��2�h���cϻ�%������'*���8��m�BL�Zb���J~���t>)d�˖Y���7mQ�t���9��!�]�+#D;�'Rr�څ�D�-���HOS귦U�8V�j -��R���w�V��cC���v<���_�w�� �5=Rɽ^�+�����
�L	&�X�z�K`��(^#���f�DE �h+hZV6�`��d�Q���l>}9���
lv����P��1�3G���˔�!��2�]vB���8i�uO��S�c T˓�a�
#�81��mW*����#ٶ5K�%w�������Z5���_����GNH� ڀO�Zd}D��"�R�ZXv�|j�lJ�ڑ� "5�h��[`H5���g��[dd�5��_�uy�PH �c|���֦�Y�O.D�5D��:��9��Y��.��TQ#�t
������
�h|\�6l���
SN�N��;��U����U��f�,�r�-���6��_]� MI�	��{
J״vu�_Z��cf}<�gwH��Y�x)���4�R#A�wV)���xu~ps)I>9g�:_�4�z��z|���|�c+,a {$�n(�y��������y�����tݢd���ae������NX6�n �m@��3�}�u�Fqft@j�I���ե�I3\�gphO!D�`x�9O{Cm_���3�to$�f���G?�w�Gha�@��9y?��h�����x�^/Gû�c,m���eH�{MX!:��(\u��������	,�f+������ckZnl�P�pXG�^҆������(p���V�cqgO]��+����!F���	]}E(���ȫ�|�Q��K �-[ތ�Un���F���
���ޓ�ht�t*�
�Pk���~a14���j�\\&� �\��P�Ƞ�x�s�֌V���[��j��!7�MLH�0�Da�G�/�%�w*�%$v���W(ݔ�}P:m�5"O�#��WD	k��i��F��OҼP*�`<hNya�{��*Ql����l�.����5t%k��8���o@k�r��&"K�7"�Ԙ����H��!��g
RɌE�������0�����[E���4^����i�f��ow�����S�,�3�6�[���4�a�:�Ν�V��_C�L�.	�v.+ţ�4�{rي���Z����οBn�3[��P)[�&�)@�Zï�B���|+u���E�ͅ�2O*�L^���s��z�.RJj�`��}���!�R�)�F1���ʝ�nI�����BS+�J�iv�"��S���]s����i�+��]��	^��y���O���5>�>�}�z��>���!c�Ց� mI�&�cbք�e����ʙl�yY.Pa*�)���jm��٪�@F���?R)7f|�oS�~�)|�(8�	���I��8Q���Pwc����e�7e�a���@�V�(W^�����������i����3M���p(C�l.�ۨ�2!��M�_[Mo3+c̬/"��Fi���)�0�h��ԗ�P\����Q6�e#sb�fh���\�Lb=R��bJB��gmG�?��\�o�+$�������]�MsLt�}��SPV�{���s�	5��?����{�%�b��Y�� �v�K�4[���xvi,�U�[��kG!�X2O��A!p����Αק%h��-	�Y!�[o�|l��8 ��y��`�=��ᘮI�هj��~��
Έ��o�lWїF#�aT��R�=Q��l�.�U�K���"���Q�(p`v.�yf�kB�C�ًw�N��e˹a�!���s��CU`�U,֙��ғ�Q.���D�c�ԍY5�)B�|�i�]���u�H��L��0�"�4�`����J� �Wv�;�n�z�0�F�ĸ��ͪ��"��?)5�ֽM�&==\Z���+��p���Kf� ��*|S9��2{����ltw&��D=��)����b(^`v_>NHMO��O�o(�&�)���V�X�J�]!�4w�M!�L��z����C/�N�4���Vv��Ƌg�V?�p�8�"�!C|h���x�3�~ej@���)9X{?� ��vzCv��"
ic�;�|��<�G��#��q�zjr�.}���F��aK�[{�	x��D��� �X���r/{��^d6ê��!1u��<�-�>8!�fg���;���}-
"�^����d�	�]z�P҇w�R���kS�e�1�uľ�Y�>���Ү��f���DwjO<
Ħ�1�*Jr�����z�Z�1��EqJ��vX��\Ч��q�hA����"v��it��
x�*��5Y����1����H��;�b9��t�*�T�7��Cx�yv>ÿ*�u���V,RL憾}��i���~d�7g�)�5#�>4�= Qu�kw�ۉA��n�'
���en���Ĳs���$T�1n�F�T|�oa�rbw:	��Cw�(�`�����X��B��?�M,n �ūYtgD��}��n%(m��+�M�J[DL���	�Ob�J�xt��wٶ�Cj~h4r�O-7�JlM�_�<�ׂ��(5-�t }��sԎPA ��u�׋	���ꮃ�b�?�!���s?���`7��3L������r T�T$!cVР6��ߜ�FrU#{?�_�l��%����f}k�K'_��V�#�P�,ڭÆ�;H^W�6�h��!��g����MN���� �%x
��)�|�j�T���=��n���kro�0���֌�qXU��(�.e1��a�]˹�;Y�(�yl�@t��kr�1����dM<�~�ǻDJԙ�Wo��3�o��¸���B����w�6F�p3���l�'�L�-Эh
.�ܘ�%�n/�v|��8�(7�x���[W�}�u��S�