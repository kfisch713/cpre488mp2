XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�:w�?��?ܔ5Y�A�=�'Q����PN��f}����X�P��_3U���9!y���<�	/n-	�z�uMP,�O	 V>O�w�$~�;�����,���R"����pAԘ"� ��|������1���rY��=%[�t��F���� ��ʣ�D/��5^��>�X�Bp��JBh�� ��y(>��W��/��Ir�ۀt2��3�Vm0˧�x$ص�r@�+v �Ut\��H�[9��/�*U�Q!��/q(�&!Z���pJ~�?{�v��d9R�J�����$�6����z�!E��7"�H��E��4���%m댁&D�(Ŷ~�
��6��T�:��w�8@DI��Ώ�l@n�F
�`f.B�����¿͞�{C��{��F��j��KRb�n���nvҁU~����j7�ǪAB�8���� ;y�ER��@��ݨ�$E0:gX9�|��p��T+�Z�iHf�i����5|˺&J�$Z���T��k�vF��Pq�1���~�̯J����A��؝=#����z�)�5�ݶ�+
WY�h����͢�y�O�u$�R����۠*�;M�M���o}�LH�-�F_qw��ET��<����}�0���I���<�Ƃ���K��MX�-�M��uQ�Ċ���B���x��xڃ1���?��`tu��N	���؜�Bb����5 �r�t]�̶ev~c�6��۞�,(��zY��xԌ��4���]ӗ�&��x��Wm�XlxVHYEB    fa00    2a40uܰ��:f��<������3�f;J��q~_��%�R�U����-A�yx�:�=�˹u6�+z����08�`��x^��}ڿ��,���NF��f���p6�<t�x㴟+�P�TN iB���L�1]3��_o��N] �VMd�u�"3�8�|o����� 8�3)�Q�@. "+G�ފ(/j[ۚ��@�Ҳ�jX�O�^Y�F������!��$��(�w�\�J�b�R�4�7�����cc�T�LƄ�B�:ʒ��N��Q���<���G˜�i�����ßo����Lgkq$U|�EW�S2$�������I7�(���-X~�3�{�e����sN��*��ک�tc�sG8��8��/�#Я^a�B���A��P�M��:G��{n��E���}���Y�vAn�y�+u�G}'�zb�����v������3����'2�|:=��! �w�g�_zW�`�Kn�`��E.`H��2��L�� �Q��7�At���.fp'��4F�F���m�T� ��s�c`��q�9�U���딸C�-D�-	Λ0g��c����S��Z�b:���S���oȎ�O�.�1늪����^�NS��,��U�X获�BK9����i��jfbG�~��/�k~X��z�\�J��z1О[
D�~od/�kg�4T������ K�.���5�u�x�$�'�q>�L������H��cuWm2y��i�@k�qA�P<����m�ǜ���ng�R"Z�{_��?�����}��Yn� ��E�6�C�:���M���$�(����ބn��!�Zp:�{8�����6�`)i�P9I�Zi�"�hĢiG
�~�¹�2�� dv��z��\b'Y#���|�	'_E�6C����Z�}/}I��R�(���΢�]4}`h��Y"��T��UU��Rj�c���2�s ���%����W��Q\0M����Pt��-g!n��*��ȱ��Ϳ����$�n��d�ωo�L���*owL�Xz�m���j<i Rbc�v��f�����&�����#uȉ�/w���a�`IF��5�x�#ی�U��)-�L�J�RI���q��8@L��e�
��[��~Q��c^��7ҪF�[St}J�nf����i�[-Ք���>�����}r��X�B���l�q���,��3�葠AT�=��{l0�U�QD|+5[.��x�/&hz��$w�n�4
+��ЅB�@[�s���X����R�n�����2��zR
!n���ݢ������&�P#�A)T0������T6��g@��������b��E���qc,$o��$�ĀO���&3 9+�)T���X5�+h�,�KHTj�уn����u~
@��1�7 O�ck��؍V�s�'�6���R��Q��iXs�oW&�$S�a�ݝ����f$B��'~���^�	u�DfGr�t����(�
�j����I�T&�m�O['����^� qj��3/���A�fr;#���M�Ùg`
�f9�>ad�n��M���_5�t��b�֘��n����~?:Nwq���'*.�_=ë��Ɩ�W:���)M4?��2@dK,���4�E�Eo��)�r�
�:K��d���̝_{닮��=�d�OL�l1�e�p�쯙+Z[�H��9�AXcڣ �JX'�L��w��"�5��/P�i�T�'�ZĊ��<<��!(�&���|���?P_�&�q�����/��|v��+��H�!C;�"���
t"u��%�җc|�"���c�"e�	E$0���e�^ұb(L������ڏ0	b��z唏�o^Y���4�	��B����i&Ϛ�Hu���W�z�J �T��k8��R�y Phش�.�F���� X�a�R,��I�%"�Ԝ�z�D��������{���7��P����"I�ֳb����aq�X� zʼ�0�E��Y��
ץ�ۗ�U!x�=Zx��F��o�C����ńެ��x����¸Z�PġL�E`����&���aZ���.݅���L�'��+�p�1=S��I���4j�����6O>l���.neU��qز퇢��bV�v�s| tN�Bꝷ����D` �u�J��g�GK%}<�PU�v�;J�G��h�����b�����7>�:�k1�p�8�X\y���ߟe�'��@W@b�2��>&�u�^�..�� U����"yc�Q`.P�����SaE��9,�.�QX����i6����|�>M�������[�4ڒ=ϫ~n�����9���4>�j#}�O����ݺ�� /����`���e85-�H�YDa�y6������=�4t�Ȱ[��;,��]�dWߴ�x/j�Z�s��mM\�͹�7"�����"��P8�#�U��WW����n*n���]���ѣ-4�~_���)�HUݠ��ܘ��Y�� ����ب�������f
�{>�*kݡ�}I�ŧ�\ Q{&?���ۮ:� `�]G�_�p�3h��>��¨1��jU���q=�#8�c�Z�V|k�>�^������ku"A���&Y���� v-�*��dudM{�UbA�@�/��~X!��Wb���{[���@L��d�"��X7:��Kv�u��S�w�E���Xެoe�5S�\/�2#�l`�^R%�ͤ2|�_!4���
Wڥ��5�a>z�
�����b�m�/⼠ƺ/Xۧ"��z%ɷۋ ����@$d�!_H�6����@��/��G������&#�r����+�+��\Yh-#��q�w�z'��{<�o�"��o���9Sj�9��b��Qx�k��Q�I,`������*d�A��Xs��Z��]����d�jO�I����Y�ͼ����)�SH�ΟOhC+X+��TJ>�f��Q�)��*Ie�� v<���^����I��w0��q$�:8a��E�zg6�o�,��s8YN���qC�d��e��h׏�R8 �4����+R�<*�jG���4��ZT��(��9�����:��p�Yl�bWkw�t,(sq���7}G񸍬E+�K�^Y��a'���/�p����pK���G���XD��_M��(�'�bft'_��tٿ�'�Ƀ
b�a���x-��MKT�*:!�#kL���-�p� ����)��fAą�a���r2��q5�LOj��>���aί"9k�����8h�:�� Ɋ;���%J����e�m�[pu���my(䵲���5dl��1�k�䴌:2uOo�!��C;�;���P��Ե�"���;qr��܊<�+��F��\��g|S^܈a��''���D������K�M�����*�KҊ|��n�(�G��G9t��V�u�W<	�s�a"ӫ1���o6GQƼ��|�βy���!�^̘p��g��^@`�C�t�����9�i�H��q�S-u���.� 2I��V�~I�z���"�KUӠ�Ɏ��S�K�֑����[O�
f�kKT�+�@ �u��s���pgz0�?D	���mKX�W� ����ΐ-���{afT{�c�$-��sN�{�+(Wz��%,�<@��Mތpp�r�� ��?�b��M8۫]��tSqFC��h�Fn�B��̝��⥯ܨm�q`l�7TE���4�|C]�KgK	l�L��qLY3�B�3�����r�XG��}�a���pP��jLA�Nx?��psuN�츏��D���'�����´\i���R�j�#�QG�h�)���f�?%�f����ݠ�)�L21P���W�~F
A8/�@&�����=_��y�����9�*뷨�V�ދ!��Q7T��VCp�(
,Ɓ�������\i�m|^����n4SCO��w*�T���R�(]������ڇ���[Ւ��4ӯ��>Vq��7$�⃯5Y����d��י�ց���yO�Q{�k�"Q
�d򲴐m&Tߧ��7��;�����G�(l�i�.�oB����=0�7b�� ��Q��~]� V��Z����@A;Q�tg���Ժ祩��;�*��n �o7�j�D6������s�j&H������2]͝��2m�+xq�VJa�� f�_{�<������-7�2#8X����ӭ��� *��[b&��`��Q��I�%*!T�Մ�g�I'>�V�������к��}����q���;<���E��<���E�]�U�d�{�ct�)�tm�;.��L��X���9n���dQ�Ց��Y,V�&�6p�f� Qg�y��;��ٛs��w�Y�W;|��C�!.�����CQ���9tI�kƜ�i�o} �*�wh'�V���������������:f{��|mm�b�41�&k�����]�eV;A��`�;x,#B]5��	�i��~)&ᒼa:d(�WDQ�G��I���}p(�G�e�-����\�nB��R��"n��qɅ����9n��ŷ�j� Cx!��i��-��Jż@. bOv3de����V ��[�ſy��[-����G�rդj9y��iٸ�yݬ�O�1
o{Y��i����ܲ�d`���8Ҍr�JT���te~�洒r����z�i��ΦKhl��1=�싻�ᾈ�f�8�7�{�R���K?u�*�sF�G�Wv�u��o`��]�9�Hp�E�Z���q�����>��:I�+��K3�j8@��s���ֵ`�RQx�~n\[E{Pk����dς�2�a��5��w�Oj��X��/�5��f)hC�$�-�����I��\��yO0f\٫`50�b;�N�1Ǹ`�1�����)��#+���q�p�3�^�e%��|1>�d��R�x����7<�@Ȋ1�1����jk"�ZY(~��.�쏡��EI�S��dT�@#����I3��i��5Tk�bO(���L��q��ʀ�ߧq�q���H�����``��U!��<��PY�4g�}x����J/Y��{w��LB	����[�n�� E�PV�?n�{j� *�)�;�*K(Z\���"�������E�ha�忒�����J�t���%g���@��`8ܺ�>��?r������ɨ17��c��;-����݂&��z��օ�e];�S��.h9�Fn��q��M7S��~��5��������E��"[��*����ʯ�_^l��^�.��t7b��Y���~ �#A�(�0~а��e��&H|��-g.M��7��9tˡ��,Δ��d�-װ��A���rx_�sC�cO�I��m�����B�>��1�![Ca��,PX���2�!+j1e[���t����fu�'�����p�!���fc�A���8J�L�HMN�t6~rБVOx&��́\W�pd���M.=V���:�A�$� ��ay��S�|}sv�5!`)G��/�DLS���H0w+"����A�^dCÑ�}�.v��eJ��B5���/��H0�N2���-�>�M�z~�������"S�&�4?������D(<J�]\\�x{{*#P�AS��_�l�Q1���[�&3����WmN�NӇE��g�d�����C[����{E���ۄYV5D0�W4БLT��Z�q�-g�G8�f�v��>,Ei1���M���M�ۥ��7l-\G�l��}�I�^)��\�׽���4e�1jǹ��B ���r�۱i>\@��_���5Ⱦ��O�%��P��+�]�#�wѳMx��Ʋ���s�5#/h��J���0pfZ����ʬ�Iku�8��0e�y&o[T���k�+V�!\��ʕ�|T���z���LP��MLu�O���Z���6���!M�:�ɦ���'�����B���@��Ţ�+�7B�$c%#�Z+ HM�K��� �:�z~P��D� Jbu���V9��X7��R�I���I�
����?��[
��[?�@\=u�8�����O��F.5�u8��gE>>����0p��K���ْ	^���k��b� >Dԡ(����"en�����:O��_��s�p�/�Qn^����u��"��"I�U�9����
;z�[���4�k�K�|)���;���=&T���
�ċx2�d�1!IԲ�����!���<�,?x�����b�6��Z�!�Y�;e���?m^�
f ���h�Djӄ��+�ߝ] 6��t�w��IzHC�Ҭ��O��G�]���!�g������A po{g���� ����l�t�S_s(��P�z�s�[���F��[o�rb����If��	8���H5��~w��Q�+�7�AZc�BP��Zo���Sw׷z�),�%q@�)�M�����N�ન�Bx�F^(UT�L�c��lUZ)<�9C]�^֨�ԓ2��j�I�;̶s��H$���A!�Ur����d��Q8g3ٮN�ojtp�Q��$XQB�M��K���3�w�r��=�`�nQ��rItj�y7݄��|�C��
"g���P۰��S�_ʓ�%ςL��d6w��Z%��bF�>r�+�~����`k��4����,!" �l1�����s�h�k��'`7���d>�o�ȈZ�*�%舜{���S�ͺ&FV�Ǟ��m�YcRC��+}�ˢ󻲅�/#�� N-Q�I��i|�g �2����b�r$n���	US�"��<�B
�ɱ�����U�P�3_<:s��X{�|٫���Y}VN:�Ѕ�
���V'(	����ZED���r.dx�����԰	���{��|UԨ?�Z������]p��@(`��ש�&� �Z�E�/�a�%W���l�*3���.$}�\�}G����N
X�x�S;���1�e?�H|i�����na���R�������r�H��,��
y��.;�L�g� ��3`"�K�ɌUH�W���&4]&�g���= 0u�i\��ȫϘ.,����{`��ٔ/�cU|o>c<����e%�`�4����AS?v�.n-R��mbG��+����A~���5�������|4|��	�w�X;�w%Y�Hx=߰����MY̧�0�c��)4%����١�->-��8�D�fR�9������M��pMC���9"��v����|%�Z!Ƿr�^|U��7�fCo��MԞ�Ǐ�pz`]A gIߗ�}L~�j<�y������&:�~�m'�Ef`0�gA-GD�{�%�)�z���Úֹ����E�<��O�B0|N`*�t7�c�7u%�!M';Ǻ�_�c���c7�;�}Yg�A����D�����C\eA�)C<�n
�����R�u_4�����z�Ύ~�f���o�14r��g���q	G�9( ��G�hן�`�}xU�C]-�����JcQ���TLt���Zl��s�7N�ܠ�q?�����)�~gγ�q<��Q����~��4�O��z2�U<�$k�Y�wnV��2���Vq�9�%|^�/!�oR["�M�E	��˵��5[}<C5��6�\&�&Ւ�lK�RS�	��I�w�V&1*Od�W���I���`��p>������ò���,I�}5y�aZ��c﷋Kq%�p�������!=[1U$��Ez[���`)�_�3�t���2�Z�s}�9��c�>��{�%�a�,G?Ś�~rK�u����38�y���:��Ѣ�fZ���ggX}&c�6�+s���v0�^M�D�e�aP
CMX�9�����Tm'9#�b�4lQ�!�ˤ4���=�������N���1]�耴�� �X��}�Zʿl0�����3skV�Ԧ�)��P>�G�.��waTSzʱ��dS���w"�{_��"_�uc�޼�2�|L��~k�Y���W��6!?�'9����'�3���'g��L<Hk�ߗ4[� NUk�8t���
\�����\��/��F��g��C(Y(���>��
_RX���,k����W����֯�a�	��r����!���P�[���roy�>=P���ʌ�!���A��f��vQEp|��J[�6��<_��yf�Z��TZW����?�h��L�q�sBZ���x���/���.�'�����3@󾳋������H�����N���8��)�һxN�\W��z��3w��aȽ�qF�u��>���V$��(0_~�33�y�� n�Q��D^�<Q�@>����~���b���VΝe�|X/�?���:�Ve�e��_ �տ ��ܪw�D!7�4�Ϲ�X�rs{p�#�]T���jԽ��:�"��_*n�wW�1@k�s��v�8r&`�*j���W �h��p������@��2�?ׯ�ƶ<���3H �Sm�o�}��p����%a"�R��`�X�S���=3��`��d�/����_M�C�:#S��$��C��3:�єc�,?���C�2g�'��*��e��t,U�j_�b�U��(��͎�I�!��Ie�H�m�z�����'�[��I� �o��������Z�	[�����O���o)^S���s��S�/�q���+
��X���Ǆ�6ې�r,Y�f�
��A�n��V����������ăȺ8�2�����Y+�/�OgA��ـ������n����m���,ʰ.d�t�:5��I����<E3&
b��֬$�+���Gy?�#K�g��q��B&��w'@����n��>���fe���6�:q��>�p��*���hۤ8!����<@��7�44�9�)o[��D��Z �6↔2�ըvS̀r�ϡ\r��u�u��1�!�%��a�	�BuF T�p�&
���N*����,W��M��%v6��e!���t��%�����N�nO�C�I�&@zX�q��f~<ݳ��!�'#�?L�A"y
�m�e�{!QF��2�֑��c+�$'t�Z+��F�E�c|U��=?����0��?8����2*q�wY��с��M�fV�c�R�6�@�2-þ�Ҩ'��.ڕ�a�*�a�$W^�\��mLd}c]�o'Xm��Sy�d�L�)�k����7�/��� 5 |��#�%E:���Z��W�n_�.u��}����Y���(���y�b��KL��2xFO��	'��z������P�	�Hƪ0*�>Ҵh_����(��>(!�\k�}i�p,g�)"^��u��Ź�W�T������X'��NW�}A+��q&_qq(V�$j���I��[�R��>1���U:{I�ε<:S�OJ�X,G�n4��d�"�4o���[B��/����XA�J=�j#%�l��b+~��q�^���..��}�:Q�%!_�$p�w�����	A�`�n;��V��Z�y�,tE0��]�e��ş��N�j{YX�֊�]�]hD�H(�W�@6���h#JtZ9$�ؙ{�D���ہ���?�a;�S-z8Lԁ�'�t���瘘!��c�ɪ���Z\	�m��K �[b��I�p��jP�.�U{���ڈǪ�@E{~q������-Ȥ_����T���&T�U>����3Ξ@a齟<$��I'��
©�1[�ɑ��[�c��莣����������������<N��I�x5j�	�Cc(��q���'����:Z�6�9��J��>���"�/x��Y[+��,�33����W��f��#�d�Xm#Ч�G�$����z�΀��)�T�gpY2���b���e��)�J�* sAM{���3B7W�c�1c�88�[�-�.��gf�(ή��jÁ��F��5�@�5P�Ee�~��g�v7��x���M0m�g�||Kd� ���`��H�?��[��:F��/r5��Ai!�@����JRP�$���4�x������	�L�=V�X�5{�:ӑ0��u$���z]1�K��i�B�#(���s�3u�b0�����X�r�>J���|��E�6Lp�8��Lh������y��2�i�/vEU�gs����M�Ƣ
�*&nmn�0]��3V�DQ�΀�_��,��ctD��P.7��N~��}��"��"�z�6[�V��7�$,Oޒ �](֞��(PxU7Az_�l�Yc�,i*`����p��ĸ�;�b� �ob�"����%�~-��x	��m-��`������W) Yk��|�mC�����b�<���g��?���z>޳b���tt�ҙ7N& Ǎ�we�lLir�f��eiJB��_�y3���^#R���v��;��7I��8<� �=t�{�.R��qK��d0
\�js�i����F�!��9�Ü�r�4#�ds��Ki��մ<�g��B�*�ԅ7�;��K�����a�
�~�RkT�� �~,0��֢ă����ϙ��[J�]�jLy�fz��m�ON~rhn�]�M�n���wH�l*��z����7����l�	��9V��N�K�N<{%F�.�fږP�F��Ӟ���t���x~����''.���<Y7x�H� P�>v�R�n�=�Z���M BVgFD�R��0<B4}@ݬ�6sb;�^�$i��gVT5a�̤{аi�0bڛ�F�Z��������t#m,rt$[��G�ΊP+ػ���h\��o��8��bO9ۏ��1 _���SG�1�����������`����{���px2:a���X�%������&
������KVaW�XlxVHYEB    fa00     8e0O�"���V��S�^�݋���Ʌ?�ʅ�@�s-�ƿ�.�-(7ckU�c-��<H��_�F�h�KsvY��!L#<�}��B&�n���O�o{�-�{L%�����ە��B��On�?��| Y�ݱd}	eЍR�V��xf�3��G�.R�J߷�q�̇}�=ĘQ�!� `Ȫ��.c6�v�-F�r���|3���^��lj+=,y�-ay^��WC ���aװM����Za��'�i6��
��-y@�
�#9X�ҞD~/�����i:(�q�6gٿ<)g�T�:�Q��1�ͳ:�Wϟ������:��xf3�6REl�m,�-�SN���(O��@"�V��xƦ׭hg�f���#>/�^?$�$~�5IbTc�S�w�64��J�`���Q�m ��s�K��;�I��'�Nnt�a�Ʋ��-�!��cA��։�����4}[O� ��:>���>y�G��$������!��7��EFğ���Lm����o��v������g�ly�o���/~���V��r���6�9��-||�*�����̧͞�D�H��J� ��m���-�@hf3/������t�I��$�e�0��E�A�sZD)v?ȯ�©��\��A�y�mʩ�y��?j<.��Q;4IR_���I���s��F�mt�hQ�rl��Q��/~c�*�Vڛ����$rb�.�f ��1�<�F(mR뤯��2��*�X"�ߋ�5K�w��~Y4�o췰�J��./I_���M*R�id$kPiG�B�.�"o Y�5�rD�o��t.1��D�^n��#FĿ�WfֱF�#Y� 4�D�h.����x�@ak�M���@aY��9T �pb�a�N<Ó2A��Ip�rR@��q�����j<��|�M�4��W�Z���8�J^�^�*;�8�����٢ܿ�	qn�5��c"d���w�V�#Z��v���MɦЈ4���Y���e�¢�w� $fז���"����m$�b�cd�1G@Ga���Gt��=X��RN�p��T�>*�Ҩ� �����6Q�������v�,�P�ad��}��7i��Otw�\'�����wA�Xp�q��j�r1g�J�$Ș�L������2º'��{x�o�GQ^����I� �16��]z�Y҄�;��~-��d
L�_�	��b�6�.��b#�փ?�A���¬s��"g9�ۛ�4�Ϯ�뤋����;��Q�����|l(p�R���3�7��WK�nzɂ1�V�Ų;����I�j�+B� �r�{�2 f^�xv@����0H�w�2B1�<E��h{��p�_􆌆�k���r�3�?ޞG�1�H�mD�7���-=�m�l$Sm�|��n�c,G�a.G�H�%��˖@�HX/K����L���KD�c0
�����M��8=ެ���B�|�n���ӊ�o+��&��G�P��/ˌ��B�+J+��<���g>o��
�]����6QE�t;�{L��cչ����,�m:Pt6�)�1k{�Eo��f����@��4���kP�<Ak���ү5r�CP�y^��!eY��@t�{#�.�Yb�(��� ��ί�P5�ɉ<����E��طC3#iV{��
�	]�¦��#(J��%T�I���4����d��w�}�j�`p_^?�-
'+�X"xѽ�,���x��Ϣ�e Rl)�%VȺS�H3����Kh���(¨�9hO��n%�<�����)���T=r�,q���M��̧�i�4��7�aq&�A���!�}M�Qg�K/ke�7�ߕ(�%c�H��%��7�����t��$"�82Y�9��9���������P��GȜ�=j�"�ƚ�ĝ��[��x'�n����
ɍ��S�q���e���v���_�.��8n� Z��TĲt�)��K�O#��.���B�7����1��;t�������Sl��Y;6K,HR����\K�<ӂQ��#���9�L��]��h�=C�B�{O8���u��xB�%p��6���
�ee���s����d\}����^�Q��.��!��6�7Dr�?��}q8>Q�G��7��YP��z�ߓ7���:vQz��I�������X�^|�O-c�����8��N�����NбD&85]��x���
�o���k���wGC%��\mt�l����
L�s��$��i,���Atzhj|dT�HZFB}�������0>ck�͸X�u�;����UXlxVHYEB    fa00    11102[M�OT�����A7��Q��ˉI������~HlT�#�P��}c��kh/���+c
�v��j��i���3�s�f�;�ڭG �ig�l=��֠���y�v�m�f�����OP9ccԇ��J�0X|{�����:La*��
ژp�*_�P��;{8��ئ~\'աZ��"�|�̸�����Jv����p���TX����WGX.��@]��%�㏼2a�F�簀��]��)��
{\CQ��pg;�+s_|���c���rs�Z�:�>�+�[OF�M��&
�2�y`��Z~��M&�dyV_+J�����Q꾮��К9rv���;��Պ�te
���ŊV����3�td�=iGV�k���5�ܴk}�؈����x�����V U)����s���a����5ѾV�~mC�.�Ŷ�j-�+!p�9(jZ�h����4&�l��-If!!t��0��ZG߻��<\�9��>׽U@b8����H�/�� ���F�ko�~��9t�ԟ|�Lz=�m�	�5�6�:��}�{��;�m���Zq)5R�Wr��Owt:�$\�=d)$Ng/��?m�����1QG\8�R�q�`�<R�,�������|i�ɄA��`�;�����Q� @���g�.�j¾)�nC1�LP� R˿�}���T@<8T��+�&Qy�P���>���<�|��; b��ʅ��[�u{��s�1i�{��밺_9�-^o�mrȧ
�EoCBC��B`��Z\$�Ύ��a}�j��W����	��֌'����,e�?	1C��x[n/wCՈ�5�U�y��йH&FL�T;ދ��01����7�|D�}�zB����x�p�2���ܛ����/�ה�1]HN��'��9$%	�\�ԁA(�K�L�ص9L�2� ��\ꗶ+}�]bd3�C�L�U����~;"�.bo`�5E$pN�� �S
��l_½�)Ԇ����_j��Y]2\�^�����LM���J���{���9�f+��Y�_�ձQi׸����c��QSl�:ʽ��@�i���O]��.n����ʜ*���͞y�Tt]�J�X�'��E9��d�4[�jr�r(��{2�W񦝤6��T.���ɛg��e�7�q��9�*�nϮ�#�"��=~��̑��/�(�Mu��mRj!��^(�V��k&a�=�����#߼5�C�fU�>�L� ���8�ۀ9D�V�� ����ez�	g�|<�_��?���w�ڊ���P�|jx@iP`~gr��}<�i�oq�@ue#�~L'�<��N.SP�J�C���7}�u������`\V��}�}�3{�����H��~rܣ^����	G�����g��y�eX'ť�<���B����n�ʮ,���ҭ����
�����[�d�:�|_�7>�MSP0�g?����r�!����	�T!S�\0�Zn=���u�����?�'^BHsۛ���n��jK/����	݉�*�Ͼ�V^E�-"UJ&�k2��1��X,���m,6n�	C�P�w�]�+C��a�.��][H�@T���,�aÚ~�.P���gR�t-F�"����=��u�p�8���I+t��/;7'�D+��3p<^jo�FOT�˗�uqd1�^Y�z;���U�7�<rݔ�O�1G�E��O�i��k�$dcZ#��q�o�K&"]�Z ��޹{�i(�F��=&u֍N�`�%���sOfc�
������2Y0wPH��f���) �%���t�� ��+��_����}U�F����͔	�n�!I^�Ò�1�r���-2: l���Y/�5�E5��,	  �/h�gG�$n���+n�r���kp��6�����jp'�������1�
7�J&�50�۷��$�(�z#�S���Dи���r�35��*��8�M���ܧ�����Sn�������)���f ����}��3q����-u�~+1���_�w��@�-�-c�����3���F��ӀIyA]kD��\���cWPLx�����p�Z�!*J:�c|�1
 ��b��ep�����<�(s*�N[}ғĖ(0�-{�>���{��k��Aso���YT$ pR�	D?�$����� Rķ��R���n�b��*�G҇.���N+>v�K��4�+��ֶ_��"��*���Lσ�W�i����M���D����:^�8�%��l}��|�^�5L3XcF�'4M2I�'�@�->a�"ڟg�%^�@��GѤ5�����/�J��	�e�/��Q�}���ŀ凊h�����<�~;�H��R����CX=�2T�5�B���ot��hm/��Y
 �uO�J+�Cܼ����Gid�?��	��)�EJ���V@�X�V�A�8�=�ǅ�k���Y�����ݦ��&6R%Z�ꖜL`�!�=�����<m��ω��s�i]�_�v���A�K9�/�R`�6o��&�A=�����Tt������V����.�#@8ǌ���'�$���o��r)���n���9jB���&��2ø���O��J
8�o{ @��JʳhQ�l��@�Af�-1��^9J��_�Fo)�U���B[���'��`H��ã@D~��*)�(%r�W�ޞ��5JH�	§k����_jI��t4�����m�ac��2g$�o�OD�^S�hy;{5b��C:Ψ�j��r�Zl~�i�e���t�/?6��L=4�8��6&F��Z�:��Zl{�6�&i��}
m�v��u~!��:M�My����J����>r����}s>]��.ZΧ?P
P����V�[ڊ��ы\���M�s���ӶW}�J����d��V�TJ��C��T)�Db��e�E7���3_�
L�"{N�/u[M�ka�QlE��K�x�ɕ�Ӂ
�I��8�} ��0	�3�}���S�6Tl}wJ�`R*��*DB�/2
�&@��g���:t�@�g�H�v텶���R'hW�-!�$61��i��
���rR��7 �$-+�إ����p���
�ب�.0�
`�H
��]��Q���!�['����x;-LLܤF�m{��.��L[�"S	T|a����|}B,�4���l�+�v�@�Nx@^��3���9Ej4�W�)iBg�Ͳ��=�v���ދɐ]�[_k�(9�����	YDX]��ߴP�S���qV(l�c��ߠ�`���7�Z��G3�轩�����ע/�1T9V�UU�OnL��\�2�j��T�'�R��K�S瀭�A�;��L��ի�g�Զ�E�ghd[�VF�>T�ϐ�TͲM��l[�� �a�+�0�����I�pWd~�� �ŕQ��3U�Aa��[�}�+׹{�(�1�D<��Ϥv���?���r�+o=�p��"�*�D���x�P���&�kM<y�R��b�$l�A~�UFo�9�K�C�ݸ�	#e�&,臓�;[mn4��y[]0�'�0�V�&DF ����1��cz&�mo�ViC3Ʀ't�Z��=-{��[!����>�mH���5�/XJ�r��sdW��
���8�X��?�a�i�	y�(hj��`U�:�~TI���'!����N�O�Dx�X6S�Z�g:��ЬW���(J����5|����*�� �$�d����,��6���K6*;�{�4Yw�q_�9����2�;���L\�8=�;��j#);���\N��Z��aQ��*�($�e�O[��dfŷw<�*��'��Rps#��C6���e��ێ�=}���8!
#{bRح���a2� X9p���6�'�+�'d���R��D3p)2��Ρ���0����e~F�oc;,92V0��k���d�ȱm2=�Z�^o����¢�+}�!K�`S�V����8w��ZV*��c�ׁdM�!s���fcd�fڜrS���tJfB�/4�S��w�|秥���C ӑi'�m��BR�FMf}��OCa��CN��K�ed��Л�}�.%~��۝�'%��>y=�:Û#�*�S���\t�{��-�~L$W�`�o�j@�#Xv~�1�h�.� e���΀P�[��||���;J��jU����B�U��q���S���YgA~ �Q�� Þ��ض!�$�V��vS�yF�1��h�ݻ��^���'g�ۺp�[���V��KMB�p���3�|��<x�|)��C��$���\!��R�Ģ�b����Ը<�Kgc�9�Ф*ƘT���YO����չ�ľO5�����tv6KE���J�d��E� ��-�/X�+Ζ�y�p.DlMT�+XlxVHYEB    fa00     ca0o�Q��
P{v�UG`4z����нO��2�֯�<���Qف�+��F�a9w�j:�q��h}�Ts��茔	�2%�=�,f���<7���$��&�k��.��^e�vC�эԲ�I�t&'f4G'ۤ������<~EB�+tHʥ���|��BT�0����6"̷��/?�8�I|h�����ܞ�D0�'��1�Hg�,��^��Ԛ�N_���Cj%�(j���f���������¾�_�gr ��Z�^�X�m��q��A��P0N���H[y�|�&��pБ��y!�j��������);��H�~��l�j[ihX:��9$�=��0�ֲ���},��I�J:�Y�ע(8���JU���%T��B�uNt>�����k*DM]�ѷB�"f7#�v�"�V�g����`��ZX��Љ��g%�Sm��Uu�)�5�!W!iQ��O�WȚ�ÁKCQɷ��8^��~�:�.�X�mjF�?� Oz:� %���F�jMu�j�D�l�u<v���c���=�J��A+X�ë���ݥ�CZ���w�b�V�^Q	�'�mP3��Gy��&��>�7¢e?�����������nl<}�=^Y^D&L���<��,�C�!�ހ�F��0��*gh�;�O+���w}���P�
�v�+��#|��.��ЉyiY����G�?�Pr��Ət�x,�c� �3�"�� ƹ�UC ��zq�2c7[��Bx�&P����ͩ��yɦLXr�R)��O���j����1�$WH���h�U63���K�4& ��C�=�.1c�q�l��5��\f�FU���F{tQ��B���&�yv{#�z���#r�~�/Z_�5�;��%�*�\n:�af�/��Q��l�*Tlu���9�)�+��B�6�����_�n���]H@k��ԁN�%jk[ѺI���Pd������|V��sz鯷c��$ �t�%���`	E�3W�d�e�6^ϝ����6��K�P��M�H5�̭�ݽB����d��;0cXĘ EP����齌�ba~�Kw1n���y�����*�E��Ȭ^���\���702ùa
��k���Fg���rMC���!ᐜsK�cG���ˁ��u�������S�U�h|�@����h~���N�1=���~�{� [������%�!o��'6Q��Ɩ���<�åő�7��mL�"��d̎C�|o���w_@��[�0�C�1`q���$Sk��#I�'D��4DI��&�[�to_�8�l�SueEl��|7�챊�� �(��@���#G+��M�(4N�cqm4�|dTS�xo+�u��2;KI}��U��T4��!8�tI�+��(�%�D�OQ�_�g^>�k��y�kPN�ԔM����ߵ;y�A���~�]�$g臧��F����x��D{�lLl���.z�7�'�o�*_�|�s&=|��tquc�^˰�%�r���b<�-J�֓�)��	<,'%u��!)��<Ջ�=`��%�pJޤ'��7��~���BY�q*54bl�[�\U�5���D�rM��w��t��r�)�EU���D;`^ȤQP�p�xSL����T'��(|��ޟ b����d�j��T�hma�{��>'.N�����?a�U��A���fw9�JK�˞HJ����z�$����I�5ܬ�ng;<���_��x6(����7Mr4�F�[l��Z��xt�J+NS� �j��M{��ơj�� YYs �D����fi��þ�\�z�*���'K����jۄ;-LQǗ���:C�"R'��^g;�t��2�����<�b��Q����L.�hPh�.6��s΅�;�Rn���6��?��m~���y��Ӆ�'<
�[�x$ :O�V�R��o���I�~xd؝�86:�����{ ��_d�ᰟ��> >U�酰����x��O���/�6��]f�*��3UA�u�W΅b:��世;J��I
��F^������/Iط���F%�s~@�˟-{3jo=L�4D��x+�X�*�i�!�YY�X
0F��A["y�6�7hh xG'�	��K���8��g��O��D1�}��' ��{�O@k�"+��ոmA�_Y��' ��p�u'F�J]㠅��QB����tV��!ڢ�Ii�ɯ�O5rFh�'����]/
`%Kh�{ʤ�̠}4�wW��]�m�T���Dl^����b�;�6\�J�z�Le���w_ ��'�����\7D�|y{��M�h�K׮��GE�e_��G:�Cy�p������<V��¢� c�Y!��U2�5�yD�l}6��O\姖/��}�p�oS=�'���6j��U2���N8�d�j#X��i�4)esb��4WFn�Q�����&���a=IS'ی���1;�)Ao5q(�K�	-�k�GE��z.M�96,���υA|#~���ݳG�:�<]n�e��/`S��?��-ڪ��<d���^y7�x����^�J<�=6��/(��`�)��c�n����Y��7%$.�r��A%�P������LD½,ڭ*r�X��h��y��aj��4��Q�{�?]|����!zâu]��U h�na*��_#�)��{���#�BC�ֽ&or�՛|y�Q�]4���	9\"��o5�H���s�{8�w'�m�0W���D�[�0=�,���n\aL��\�щ�IK��g����@~�4��j�B�ԓb:��ß8im�{Z�k�d�ֺ��-�-�YFx`C��(H~"��ɀ@>�LF��u��~t�_�K�ݝxl�[�Vve�O{��+�S��MxqNY5�ٷ	�	�Q����oP�r�ɒ��U�� Jr��l�����5C'h�&����\�* �9WB�Z�p�"�����Kp?}�LwCJ��6��Y�0��F���7�ᬕ��Y)��I���7z����%�S�ٴ��e*�=��WQ��Fa���a��c`8�D�^
��iH���گ@ŉ�~��l�C��LI�O�lgS�0l��c���I�״~� ��-��Q�����8>e��@�o��N�E�1�ܳ8�pۉ|3�
��n�1G�S��l�$/�,o�zԹ�8xȌY�U����gy��M�q�E`�ni�s����6�:*U�w|K�:d��e�!�BxUPX-Pj����<���044�%����{Z��#�踪y��L�-�Z���$�üڜ'��XlxVHYEB    fa00     3f0~��H{uH*�di60��q-+X���(�D<J��_ %�Pw��	�7m�8&�ah*;K�o;�mj��U>���3�1��j)��>b������=f-��v���󻖀�8���VQ"y8�聓�?FLg��N����g>$�|�O�Uj��8d�m��jx�R�^
��~_�Z(�f�b��"'��}�R�ic���w>.�ȥ4EA<�(��~5�����>�Q�/`��,�roR�ﱻ�Z/�����3�|�p���D��y����߇�I(J[�`j���I??�)�&��I�{�ŝQ'E�غ.JI�-�Ç�O�Z���ꇰC��=	T�|f9����q�e����Ƀ���a̞vA�-�N�(/����e!�|�.�Җ}9���z�O�@{N�}��&�1lG1����\c�Iʝ����[:�;�q�z~�NJ54��=0|u$�Ib�pc���8�|�9�2\$�� �6��(ݏO��|��eS��9PE>�^mLd9����An���O<�>��	n˥1,�1�D��Cm��/��Ș�BW*�>���ZyV��28��]��?��2���� �{������i�^:x��¬�Kl^S�p.Sʗj����ϻ�U�������!�7W�y�y-[V78�������(����Je�w�U=�cf+.S
�ه
��Ɗ�a��S�y���l%��)P+������ä@�k夏�QemO�
�;�}2�ڕP~��#$�bmV�M����	�|]��e�8�.~FY����\�����H��/�K�
HsDrȘ�~e���v�j8�1ȄU�
Į4R�(�/E�v1雐i/lk�j�=&���P�o<��	!&��5�o�e���h�˹�Umm��'��ܧg�|:-�ʟ��ˡ�S�:f>�!�7Skjr��؀]<����Mv���*1$��j�ڵ��i�7��M����S*'�΂�@�>"���+�Ha�TL�]��ǓBs5��z�,��N����I�l)&�XlxVHYEB    8096     b20��b:�jj������T�c����{k �k�7�	`@-���,�-\X����kC�_���������?���������&�7os۪���d�F��r<���s�f�y�ht�J���� �$�^���/���1��&�},����9���oLyR�|�+��%�H�H��>*��%|���g��;��-f�Ɓ�n&C�����tM�m��t^��#��IV��G��.��}Hb�,���Ê>Q-��Op����%�o��F'�c�;���K���O�E��	��
��Q�Ʋ���jZ�~�C!J�\�ǲ?�絽@&oI�(>����r`�a�o��T^C뿆��ON ���AF�9����1"��1d/��_S�Gn
3}�B�=�P�O�������T��]��{��Bvz=Β�*���N��i��(kl����9H^��wE����[9PF[�O
��1��˫������s���s�O�p�!����h�2�8�ޢu�#�&@�CI�lu��ه�y�����ܲ!,FW�+`��=��>l�ψ��
}�|L����3�����նwO��Ғ���D`���PZ�Up�P���.ާd�XA�62��m�Ҽ�
�C������v��Sӱ�+�ֽ
��[Z��i%��	Sjّ5��T7]T���R<�+H���y�P���\�a���q���w��ǀY_��v��۞Mrt�+�F�����{��U���z!�-��(��ˬLN��?O��$�[j��nM䠝5В�K��)�I�_7@�q�Jk�v9䲎D�Ƹ���t,e	@�/ļ��*np]մ��#h�ӱ[{׫M��,�Ї�e(����LZ4��t�z�i%����;��9��5fjG�#	n��Zw;�j]Z4������R����Z�K���4l�:��;n0�f\�K�o�fǆ�X�d��Y��u��mNu�[�;��{��>�w�p�h!aS� B�ӞN�O�m�NR4�q��K�l~z ��[V��؃����w��UṜ�V)����x0�����{t��P6s�>� ���lA�Ƈa��_�w6���[E�p���\4AҖ�75���Z*E��j0�X���c���������� ;�|�f������%��K�-�0x��3�2h���Ъ_��v���xy^�
X
����UY��`e������b������+���U�̞!�|�r��]���n�i�^j���Rl�����T�p���Z��Z�ĉע����vI̸����D��,����<���w��ʮ���o���bګ�v4u���é�ϫ*��-�Cؘ#I�:O�.~}���4��i�XbԪ��
V͙T�r��Y,��79З�q��Z$��
��Jg�=�8H�������>ZC`�.E����wR��<�YV�k�oڽN[�	�>��A�U1z�ұ�d�?�f1�>��ա(�����������5-A\���|�nv�� M����m!�ǉ���;ޣ���	5~�[���I������� \�(��>V5|�a�)|�gu�@�2�j]L{n�w�hǓK���s��yQ��H��F��:�����΋��S�J�K���0��P)^�n�?)�}R��VCp���6^�.� _���+�
���=D�b��c���o�r�֐�k<��h�x���-O�餆�H� �+s�C3R����]\!�YZ�o3r���F���!��|�..��A��:�ٜƀ�J�T��	.޼;� �:��o��s�e�Zכ35C���z���!�dds�?d�")i��!�:�ԙL����=�X����_r��S��/G�yr\`c���Y�l�U����5D]W�6�<c�_�*�sQ3?􋎫��ٗC�6}�ľkP�H����߯��orf"���L��%����{�.��k�+�'�?%��#��!��"�w�B�~*����@xH]T�����2q���"Jf��·�;�񃗊�(��<�1�����lr��zO�e�	��S58�-3E��a*D�l�-V���`��v��sr=s��M���K|�-]���ګM��UpQ�ʭJ�S���]0V��.�*N�v�H���f��Ɏ�a�r`	6Q
�I�>a���@���qP�`���i�AI�����F���b�$��d#�O����ep*jR}\TR~b������'s]6MU�ƌ���:7�`�����/,��e�I!���rm��P�V7's;"�}�k���01y�6��j��3z�Oo�6�\k	M�a���Ll��f�mWSd����ݽT<�^ut�N������9Ckz}L�L�t�|��_W�3Ֆ�F	���2@!pI�V�2T���w�'�^6�-����#E�P���N���f��]����sI����im<떭!���oO0�XZ8��0��fp�]8�ϾD�86~�z��m�V#	GFz�~_)���K��X����`��Y���ِ"6�0�ō�>�!�O��aa^'�1i�i���V���OFU{J��~z�T]��0O�E�`O+�����m;��Ӄ�g|��cZ��>o6���i�y�x�&m�bJf�L��.�QO�:t.%5�!9AIՅ�=j�|�&;W�~�������\�Vb%!�#Rf�j���߆��Ï͖φ��1�v�D��>4�P�=��b�˶��ǵ�7d���8y��w�wf;D�K���*�+$)����яc��c�`�28/�h�'�qN�(��}ε�nt�r�.S�1+���ڵx���T�qi��P+�hy��ٚ}mh'.:b����po2D�J�k��\7t�?g���d �W�k 4ҭ�rz�