XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%��l!�Hi�3�m�<�v'�)(o�hY9�<n�_�+�x:�.f�A�Oޏ�&��d���]t���+h�� �"}�K���2���'���e<+	T��?6Q^ ���1�=�
^�L�l���0�M�W��mSE�s'�O��~v@��l��(��n���5%nlӠt�H�)&=�P$z�W��n�"�J��8����K�~W��TG�I�.�UN����Q@_�3�6�~�c�S���B���<MSjV����[�ҕ�7'a��P�U��+�kB�nJ�Z ��.۾��ځ⩊[A�� "����n~�b:�r�^=��]��|��hJ"��a���f0JI���,b��j�L
��k��8����P0~�]�^�x��L�9�U�*�{MS��,��^����{]גjcY5t�uy�\N��0�y9��Ga��)����L�L����M �����E޲-���QD_JP;hȇ��Ih�'{��b>4�#��v�X1�=Q�k'��49�{��v��z:������[z�9���Q����R��\	*�B`��*�vO��XJ�e�/�$�a� �g�䲐V��
�zT�0������_7����n�_)�^��,�l�ݶmG)�A�=�ȏ�P�C���>�Bw+k^r�\���>��e(���C�$�]�-Q�����u�*�z6�*:���ZB�\G��x-�bT���L�͎�\[G��F�Wq����n��P���,�h���-�R�}T��,>t����_A</��=�mXlxVHYEB    da59    2e30�~Gc��|,\,X�NRXU����
��sҋX�w*�U���Z�P���Ls�#��_����'��U�*��e��uq-0	 ��uRu���sO�/����/0��4��$��ܖy�(�oTKsʲ� �z�U���/,9"kt272�}��I��I�����,J���˻L��;@������ZE���Sn��L�P�M���F�?N�0��z�1�ⅹ��=��i������OA�S���<�c�*G�F�h܅H~�]���+}�cY1�=�����@�F#�53L	��5v.Ka�I"�Φu�̅~��\?[9� ��ߟy�P��_&����|�yྈ�pV?.W��c>B��{?���u���޲���gR�H�+�f�ر�ȋ����y��Q��3�*�A~`�ǕZ��2�W݆)�vp9q��5���ӥ$�=����$�&�j�3�	k�H\B{��:;tw�L+�#A"�O�ɀ�}M7.�(�Nđ����W�5Qcw
��(LOR���оp�\O#_yv[K��"�j���R|�n-���p�@��#,�9�����[�o���C�
����l�E����/2o��Ta�)6EC��.N�����ZkFd,�)�[6V-��R�Y��i&�KB�y�:I���%��x��u|�5����ַ�����5Џ-���1{n�b�`��úZ�ـ�kZ�y��1*�B]��F먬G9Oy�@?Ô��#.
��ZpI�4�{����td��T���M~Dvk�����t>�!t���b�@����F^#�~^����ׯ^a7�ݣZfyd�('�rV�7��uRb��u7�n�U��D����ѥgg�NP�wB�OL��I����*���;)4V�9bku�yO�?EVT�O�h�ϣO�n�ⱖ�?ɪ- -"����z�dl���B4z�LwNO�����"���:{XL+����h�n�f��4�w���u���G�*P�
�/����ʸ�+�	E|��.�f{�!�R/J��Pb�VE�ϭDV�<R�
zÏP�C����7ؿ�a5f}y�C�(n@W�
ӐgJT\���Bo�X��L�z����N�k��c�ե��&|�ܖbӾ�雵�$į��T%�'7T#�Y������[A*�Hp9x@%�	�q㵆)D�A�4�A�W�4�2���N󝲚#A������Yu���Z� |�:� ԕWlg�F�$�Le���.�*����I��G8��;�HB��5�r �?�Jl�ޑzC�S�8ʍ�W%�<֬��Ր�,�F���+L鐆,9��R��'�%���4�R�+^���a�����:"TA�߆�.d,�!?�9_��EO)�2��e������O�qG�"�z��:��5���{������P:���3�6Ά��V��N���r؍���$��L:lS�TU?l�g���r~wn��/�C�)�.6m�f���T�P��Œ|D����[ �ȃ+��;���/�3�yh��f�b{�W�%5�7߽=F%O%�X�1��j�,�l�'�..9J,�'�1\�4}S�0�O1������k_x �`&�0�����	�R�WKU�8"�x��SQDc5�����GPx��mT��6���V'���:����nZ�G��vOvm���A��8�~%OYQu1�?1%X�<y��`�;�p����J���7�,c�� ��N��Y��`&��"p&8J���WM�Z�3e���N4'���] �z�)�)��x;�;��9��Փ�]� �Rxn/
?��O�z���G�Gj���	7��	��h��>��@�z��l�|�_�Q봋���Ez����d�\&�.�n(�"�i�ģɝ.���Ym>z����d+H�����Dlu3}({4��:�e&l�L7R(z�
Uk�,$�&�1�xt����!�F������*	��N�g*گ�5��L�o�}E��w@��:��N�D~��s�q�6�*���c]L׿�h�y��X{�w7�E=���,��w�y�@9��ߗ��;|r*`a�p~�7s�Ovm�i���6���Y �c����S�؇�AMG��I��ƛ�\�ڻ�S���j*�Y�e,���K�gK���_�MH�#��9���H)���@�O�����'�a��bɠe�9�(k�N�k�7vNd{�xżfts�ڐ�w�i�DA�k�%�>�,|����<)�����ɢ��5�{�q*�2��s����h�C�:!MN�I�*X H��{>������9Q�?

�� ��,��ZBhH͙���T��!�p���B]&E�Kc��iE�H����Á�����o��jiiCj���ȹ$�XB(pI��l�p�ʊ[�1#��l�`L����|�%�s�g YU�� X4���m��ȑ�r Α�n�я.G �*��R`��J��@�g��!D�.���Z��
M<�P>�B��vڛ�*��=�����e=	@�w���"$	MuX���9_���5��P����8��;�9j��=��3w��4�Y�#��V���m�ޔ�L*ǁd'��迳��O�ŵ"�V� ,���J���8�/��#�(+�t��w�7����e�S�AW�Z G/���6o�����o�ĐS&y2��ͨ�9�߽�g�ºe�)�ֽ2�9�[ƽ�����2
�(�)�ca��|:�<��_X71\�U�©0��j�>N͸4'�q�`��]��5	/@f�T��/���ZD�ωo����*a�p��$QDiGl//�V6���T�u����P
�{���&q�&�#I��
�d�`i���Q��[�`*��5�=�-悮C�34�@w�<XS���#�����bs~n�7XgF]8C=��ʶ�t\nT�PM�}�t��,��:_��`q.V��(UX��.}3�5��gη�f�*q�Sz�"_�S�?>^�;�!H\�v�9�L�{�	>D�۳��������M�;�͙�'4��9lT;@G��(�-��G�c��XSU}�&���fs�
���'W/�[A��"#yL��H)]���/��U�.�`�Z�M��U��H��؇���ֶ�m)��5���	��Mv���!x>1��0sF� ��6���$��)�QH�؅8踬x�4����k٫:�m�p�nmng��l�F��_`�l��o/k��D~���W�,��I��V�K����޻hc�U���b`����K�g$%6���Ì?s:л�&��x��G#)�\#7�T.��4?C/\��|%���`��A�����L�lI�e���-+P*+�E�0�4y"/,Qc�S#��N)�����+�w��X��kC�(��$��	M����*�i4��͵?!u�~��h�G(��`��A��=�M�oI(������u7�M�������<N��Dר��[���@5���q.�s}h%�.l� q-D���T��qU����M�o�!\Yq���
9� ������Jw�8o@�G�o��k�5ۻ"Y��5����?9U^�����K�ݴ�fo��m^��n�u'p���_�PT����<jJ�|�"�H�P�m5ї$��e=���^I��y��5�HL�ڮ��1,A�����I ?Q�i��j����q�Z�6D�?���L'=|i�Ⱥ��x��\+�5\���%���_j�\�����089��K�e�S꦳��؈���;�zQ'&�?"$e�<@~�$���)�%yjYI���FBz�8f�:��� 6=/���|z�	3��fc���=5��������$���G�P����~V��ڰ�/.p��񶼯���"G��,��*F��R��/f���j>��5 {t��}�9=G��e���V�4
�M7���;&�J��AQ��B����?F�d����8�'�R` ��W��^hPJj[޽�e5��V�ؓ@\2C!Kf�C$����0��o�,_C�;��:6�4Ԧj x�;䂑B~.��w���U����0��<����jҪn�Zݓ�ߞI*.�$f�/��H��d/�%�){�˔�z�hH~1ڕ�^�^����d���%R֥��dГW��3\�A����	���Zj�$����/Гb�'�q�A�97o+Ȼ���̓-!w�x�H.��c5p���q���*#�D')���ؔ�ę�tc3�����V���\nL9�����~���I_�P,������ ����ʶ�R�q�"<�[58�eH�z6�S�5��5���Q#oڜ^����sN�cn����ir��s_s�#�q�!�
�j�Hѿ�j���A�?\8�/��<4�i[��w>��!q�=���k�c��d}"S���" ��C�[�ݒp��ͮT�J�;�hdD�3@y'e_"��P�Q�Gʖ�/�����$iq":�9P؝eM���T�-��Z�\���z:�5�Qt+Q]>����y��ߒw�^!m�d�����7d�"�h8`�O �25�{4�R��"&�-�}���f�Z��N0B*�;c�c���@���K(k�l/|f���@m�`���A	�OD{�8����~d,a8�LxR�;q��az��qhX�e	�"����܆լi�"�����,Z����P�LŒ�+�����\$�g9�A�}�p�oޡW��?��BG�SI�R'?b��\_��0�%,=�A󶿎y�g	��0�3��cq�O��_mpl�~*gC�x��\?2oK��J��"p��,_��K���N���}pɌ��__�� �HW2����A�g���tdQ�IݛB� �A���y��
���(����[�	����d��܋)��y\��L|>�����A��O5�ؓ��H�H�N���9ș��S���As>n���Cp���K�����U�}Ȯgy�O1��=L1T#�G���؜��Px�b#�Pi,�5X���Z���zq��6D>�	����\��DB'�-r�[6mPT3e4��p�18�W�?�y��V�f������d�������������	(W,Ն�����5{)��'�����7���������-���?��+��Ax�l�9Z�11�삵�s��q^R��P�W�C��9�Ef�B�|�^c�T_έ�g�O�UA���Q������l�L�UY��]����h�XL2��j<�r>B�����B�p�O|l���A�I�0'*��gnUն�:RT���֙\����d@2�Ɠ��06AF��%��o\��g�D1-��z��5C�pI���:�˖�`��u@ˏ� V�������(��/� ��؇��qڐy2���P`+�YJ�_*�HD<�t-�o���cr�Q�2ڀV�>G
r��殀>`%!0��w�����'�� (-? 'P�r��W�Q�Ծ�-�v8G���d���z u��R	���d�(����y&H�6�^J�E ���pl�ڑǦ�Ekdl*����`h����;`�̝�������@�\;��ѓm~]:�0�W���|�"w/���r�AQ�J�lRckI^�99
[8�&	h	
���GX2z�	䶧��/�M��*űo��0����O���!�F@��
�Ik.��L��ǈdTZ�z#0C�#�����$��G>�9�o����4x������o���,,,��{X	G:8:���ߍdU��\�[�-)���]�4�� ��R�JXI�?���7"p���Cؠ�)�饺�X�}���8�#i�{HLğ�����u�'f��hN�m2I.KF��Q�%sFP;33[2Z�s9�q�cD#揧_7����*Ͷb�c[�_��������[ʉ�:r!�\�}g2+����Ӫ����u�Y�ަ��&vj��%�Q�v��>�(3��� �3�]���,|N1g���z��fǀ��6.��J��h<������=�}c��,�9��n_V��[���_ �k�s��݇�'�Y:�6jA2�`G���G+V���'�O,�K�PzT��"suP��{����OY��(�F���3�TF���׈�!.k�~`�%m�|#��E�О�ͽ��!�6=H����&���$��Ԫa���:�7���.���z�nٵq3dS�t����Z!l\��}=��w��,r��{�;@C�+�\�����T+�l��t�Gc;�)��q+�չ�@��P;��_�O�Pf�Y��"[��Aڑk$�!���s��C �J��cKk� 1U�'K
h���fi�c��a:*���Z[ L�Ư^�M���o�(�ޣj��{1�_y���h���o�����,);�%�OMrC��N�'̍=S��g��a����R &b����<ٙK��C{��<���$+x��^лZ"��6PM���df[�h�d�g�Ol�����Yj�; @��.
���C��QC>w�3��Bgy��m�s��f�_>�__��P;�)o��`���"���VEG��!�K�YU�E��Dl�b,�Z�g_$�Xn�ck��?^S]��Y�cqf\.���)�f�`'t����Z�7Z�U�P��<�Xx��'����X�,�����Eck��-6-L��{ݾ��[�k�(��	�N��1`��9mڥ���C�m�!.".���H��[" ��P�3�eZ��ug����3�ޚ�I��w�/�A�2�Q�t�0���V��Y#����� ����8�;�#L�~γn\�`A��m�z%���~���Y���5�A�� ѵ��X���Ca��?�w�KE�S<�deB]2^�T����^��+��&�X����.U ��|�4���DV��h"Hp��y�Lh�n\�	�ꌈ����I8ԥ@*��ʕ�����j� sTL��g�EZ�����#yI���T�ֱй��Ua�A�U~� ������=o�����֠�ħ�x#y����i��t��-�����՞ZYi�"9�{�Y��}.wgۣ?�63���*���iG`,����p	����H��A�`�k���!�s�k�,�|!ŧ�$	��\����Կ����R��{Դ|�g���6ǋ4{$"�ˋ޹��(�Q	_�w�8�I<�x�"̾TLk���L(�k�{�-����~)'\M��6�sI���C
����Cy��7'����4#�T$��y����Om�Ǚ{U&O��|�������8�w����l%֙�'�~ ��NK[���镃��G°B�K��t��L~*��{)�u���f�Bݻ�n�@&y��]���� ��c0�`����8$�嘀 2M��@|���
F"���p�J���xl���?g�S�zտ���j�|��y�6�.滀��	�9}JT]�l;����B��e�(�8��?��̀5��G��ڟ˩h�߹��!	e�y��I$�8j�S8���^= 8����&�7�?��6�o!�crw'�#���v+��eDO�L(��k"��y��,s�ц��-��D߸pg9o�%�k��k驉Љ�����a	��8uk�w> Q?�2�jȾ\d��Y���`�A�d��݊Ӈ7�������h{��nIYɰ�m�l�ڧ�/t�@
/3��q+q�Ї�w]a�p��q��Y�Oֻ
Q�1��T`�����o{d�"��<n��y��:h����"�����n����.s�ܫ,�F��t���+�P��3ڮ!�����,
g�Z|� E^??R�����|�;�l�9XqP�>m���8�����ۖ��b�v=�� ac}��ײw��ɾ��D\�#�������"�a�2v0��Yg��s�;z �H\pb��.��L�o
��#�B�52c�|�������I�����ń�[�L�"2�S	m��B4�c!AJ��b�8�b3~���|�!De��ԀKm1��Z��bgb���ʥ�~
 ���V� U/��|�!C�����d+N&Z���dc*�ĺ�J'�����rMj���l�2Y2e�>��j������E[Q���ny�_>Z��#�d"�nN1wv�%pO��W����B�D��~�++/��P$�0�|G����iv
���z�L�f�����>b��i9���H�v ��,�~�6C��&����������Q�����wq���*�U� 'y�7;[h�p4��&W!%csFB�t"`�`3��6���׼�Lia�T�Ӟ0�j/�kN�+t�x[��I5��9=^BK�r�<�y��r1�	]�5�b{]ku����:�����#��"�>��x���Dz$Sh���Ȍ�҂~Ӝ~15)DI�.�_���ޞ<Q�0�� 9�$�~j�KfA�n͋$��a�E��'�"���K-�����}Bh�G)�j��r�Y�3���߶'YSS]�U<<"ax��T�B���%���S4�4��T�J|ɜ��EP�"���9��Ǹb{�c$�`&^Y�`�*��`���<Y@��~{��ƿ�ScKS�k��㤇k&�Q����=$��u��{�H~ω	Vy�اy�|�U�Y���&2�q����Ay�%������i/�}e��X�߰�m82_4}�(�l�����N�^����"n�k1��sqyyݙ����v��	%�2Wܬ&�O6\�xQ#m��؜K�,1��d�6Tޚ �z�'�����X#�U����Fv�A�0��4���h�آ&��ͤ�x�@����ٰ�wK�F�|/��G2� 4�;�Y!2<�ѳ�C1�����8%42���%5���{	�A�B�7/
*幁Y Ơ���@��D�S����'����0�g��b4�Ԗ>ٯk2��߀`�����ஞ�}>����i��/������Q�S��U��b��t�^�8����f����74ҝjn)�<Y��Wu�������Q��fW{jl���hΐ̛��KN �6� ��{���&� ;hf0y�< (��P�`�7߯3:��w��Pھ��x��hW�I׀[鮜e��� �j������zC�\�i���y	���b��ӧɸv$��F�vT��Ά�N:�*�i����T@�f� �CX;�a�����2ѐ�*,�Ӭgxћ��f��2I�?�@T3V4���F�8�
���/�k�'��c��Q"dX�����2�`�������������������BT�W�Oé`.�����ǎ4������Т��֚�����������2����K�omv�M�E��9�\�ʽ.Zzx���lC�B+NK�d���B6�D���*�����3��_�s�����4.��`�۬�)��,���U�D<sERM��ȴ�^{u�aج��i}�A\�!�B�+""�X�#��`�4���W%�ɬ���gl�C�M�\�:�R���W�!����8�ѿ�TĪ�� K�/�u���AVe�^D%���ߐ�b��!ak]q��KB�>(=����W�g8:��	�8�)��O��1?EWmo�J8�6$�^�-�[�A��������@�1�`�W]9�Y>������z�΄��TW��y�y[k#��5|#JN��/hJ%�>)�1,,
�9��c,R�~�����%��u��E}g��	�g��6�������"�՚�!�#�,y�7\�"�Ց�hdJ1e��C��׷�q��(e#���?�^�GdD��3`\�W׀�Dl��0z{qG��_�a�F`CZ~�t\ْ�|�,`T�W��R237�g��cK� 5�����Q3>���*a�N��� �_��پ"�o��v=�_+�A��A��E�8��e|��{�
�7���5��o{��)sC��� �*��8��i ��bY�TlS]��5��R-�٦�|\i�,I����O=t�%���O�i�Q����/�7m��*	��e�J���E|�?↏���a,��)�}.�ֆP���X ��S�Hn�a�*�g3:�D��}��1[�t_�=d[�ݮ���$����g\��G�~�&�`�a�E�`����0{F=A�r3��vvZkQ<�Ϫ� �x}}��=�(]�X�OϿ8��
8�;�o�T�sR��mu��n"��૚bnL�t>�37MOȓ� ɡ�9����@�KG��o�h���]�~�*)Tt�i?[��/R6S��y6��f�`D�Mp��5� �e����$)�����_Gr�W�,�.���z�b�U�.L��%�8��ue����o,�@Z� @�x��m������K�3��+#v�����RU�d����#%o�g�,ˏB%d�6?�H�v��~�+̪���j�9�Ζ�����ȅ@55���滁\�%����s��;f���J�h���%z*e� ����Pxw=�2o�G�°6�0l	��e���P ��b��֖;�.ؽh��9��h�tm	��0U܃/�U�,��K�J�=�V��!�2��-��q���w���ה:���v��E<���=����BƉ���[P�Qi�@#N��4m9���(��'#�Vq�H���Gi
f��b��] "�A e)�~�?ì]��Yȿ6�m<�s�i��$��\:�Brnf\� �R8yM6�۝�I�ng���5�v�إ �4)%��B�7x߽L�L�A�Z�fek{5d�MD�J.�:a�F�OQ�K
䐷�&��QD���M�	�\��5Ag��%���v潺�(��ـI�[*�=[��Ca<!��聩�S�� rXǪ�(,փ��$��Ճ�'�l�U �U��F����~�<q@�6㪫?���jK�S��p����V�`��~�쑊�	@ly_H�Q�8����HK#[C��~7�V�lw$�Y�[n���#�5�d�Y�ST�T��!��x(� �U���vBn��`:��)�n ��)SY�D��T����`�`�_S:�h7u��{�W�����c�3�x:P����/Z�Aqdр���P�w9���q��#y~�Y�n/@�����]�њe���Y�M���A��b�v�p�̉k�I��6�Z�yCd���W�C���u���X����._)�bu�q�^
���,0}���t���Ycf�x�8��ә�
e;(گ�FHq���
\�����EW[�(��/^v.�
��r$B�@�c�ox�6 �F[L�#�%K]��є��S����<��6]se��H�B-�g�a��bTm;-٪4�(ǇTx| Uz!�%��y~�+Ԍ5N�������\���U{��(Py��6[ҟk1������؆��x��Hs�xA��� c;A���"f���)�& �=f�O˄�?������A2+�-"�9{�92#���jpmw��2ԥ�:.MѰ�>ɁYʺw�塔|�_�1h%�0.m�*S@��	:�v	$t����؟Q�6��������ǥ�-S��J�݃�f���b�$>YU�<�r�I�����d�［B���x�ȸ���F�	�GDq���P�S,�l%;���e����0YNf{�q_�����A��o#���ɂi�ZV2�]f&[�WbZ)|Ɠ�1.�F��S����׬��,����&��nbHY|�x�D����і����}Nz�rlA'=���yن�2Co�����=k~��K�BZ��bڸɏ