XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<��������������7B���-&j��]z%�fbuQuGD��풳��3kd-��0lR:?'�j��� ��`�~�9�xO%`��1N���^ot��MV�8�]�v� �I!�o�u����b�g�'Zg�@����c�J#�4��|�W~{��Vb�;/F�+�"4��L��|�����A����| �b�8z��n*����	���-��8�M�F�_��x��Yz0��g�G�F9,��F�'!8�N�
	�Qe��PE��l�r >2�����݂����n���@Q
C}L�ޕ����Àg��V̇5�����2��
HiJ0^�5d1
�9ٝn�K��H_}�1�r��J$
�s�=]�s�9P؟	�Ġ2̀���wJ累��LHy�D�v�r����(����к��	��L��p��K&z�y�A�,4��?���ܟ���n|���w��^8�0*�'M[]��lZ�A���j��˷b;����r�.o����s��j��"��$O���!�t�8���+~�oB����P��ސ��*,�ߟ�y�3�!C�9��XȮ;���l�FN�
�ЉF]y�M�hO�����"�:��Z4F ��G��:*����:�/c.7sB�d"mq�Q��M�f?���`1��
�o� ��8�R�� V��9?L?�ȅo�T����!�@f.΋UB돝39����/����f/C����5/D�.<�?��<*G�_۠��+lxȦ���0�x˙��S�.UY���Vj�XlxVHYEB    fa00    2040�(����{2}$:ҕJX��([g���VG*�+���t�[P('�+˽_�I�D�����ڽ�`�\"֩H�Q78'�1�tW�֝��jm���Y`�o>�M�	g���"lo"w1���?dy^�:��|��֭Mo�fr��' �LS=�Gy�X�i�:�C;@gk����rU�o��ʬ媪lpN�Z0�Τ�m���r[t`m{��$;/Pb��.�I��1��$**�X W��k�+2j>�]�(��a�����������μ!"I��T���x�0�q[<�%{B��sZCc|C���Ǘ,I�@�:C�"^�%8�T��X�.Z�m�ћ;j::4��������B�$�^�@��s|�h� �v�U���`2_�1�	pc���`��T{/���n��N����c�����6+�mq1�_9��~��V&X;S8��4L��A�BKa��-f�BtـШ��f�[$bD�a.����|����3H�<��g��Y
eO�!�Mf�h�,H�Ջ[�)���ƨ��U�=������6�4~%+8b/�n�J�`����������Q��hxt�N8D��E����� �y��)���#m��髸/g�(��y�3(M��u��b�ǯ�.<�v?a�ҁ���d5[���q
D=�W�ꌑ	�L|\��Y��`�||��t��۔^+z]r�Z�O:��x͊~1�h��ɤ���]X@U�
Hp_�'NMk$�����/xn��S���*�ʰ/�i%@��E���0���1wG`���L������̆7l�x�d�:��r��H�/���no�Qן�G��@��魝vL2�=*8�y��#f�>Ⱦqy޷�r�Cμ��=�{�JI�-�����h��{�i��V���yâ�mUaC��Xz�<;	!%�]c����a�}U�c��^�����(���e�|$��Zn�{�r0�'In�c7��<"��!ժ����͉������w��r��
��t�q�p����)�n���x���D`�!�ʹ�q�1��<R8������Yf�ǿ��Lƍ�55`���E�:
�rv�k_��pj��� ���;w���Hr��#�W�|��4ݎ����ju�,��Jl�j��+�9����Ct�x�a�R2��1��1�F�Ӏ�d�q\���f#V�k`.�x�E7|��	�2�3c��
�����<}2����tM&�d�DU�,���wC> �o
X�9g��
�����H�p��2j�4���n��[��M,3��^������uc�~+,��E���3�V+��^K�����l������V�c�;r�J�i�Lo������7P� �`�!->�Zt�N\����.��H?�p߶�'"�	?���*���4���'��������l���.u�S��O������."?0g�c�w�"5�=_�*��i��������{���%\#�ny֯�����wn��cK
m�NYR�C�x�Qg�?c%��l�ЕiP�X����RTudt������A�g-��.�7blL���e���`�ǘu2�^A�C8�W����V>8�3o��/N٩��\е�3���AMSX�����k���9���V����.�N��m4Xs���Λ�����4�	���ۣ�����)�oW=F�H5��=�!��H�q	iQ.̂JK��
].��a���Vw���#;);��eB�rh�ߎ��-��#��IcdfN��	^is~<�˱H�68�Y���B�J&�l�H�$
���3��qd��N�k�5��,�1"�
:\�����8NQ`n[ 	4�N�lp�Q�!_�V1I�����e�ڱ�n�Ԭ�(�_����������t+!���ȅ��yU��_�N��rٗ��0��y ƪ�Ҥ�E���IJOF�F0�YGUt��B�[)Yժa3�2t��A�@��X�pU�nD�ƶ��U��IB���D�3�k?4ĳ�NN�	j/-#wQ�C둇����{Q�c!.2�2�m2K��{��ThG�gX��~�3d�;�1�nYX�Q��zo�u=	���#tƅAH�F;�^ڜ������<fp%��ۊ6�JB41r��H�'�`k=#a��'�J������k�t�6>9���^�o${����HҕV��,dW����cC1a�!C��ٸ(<W�{S!O����OI�U~敿�Y��p�oAG�,����qfɲ��>�Mϫ}��嫲p)�F(�z��74���(F���۝��Q�����+-d���A��U[鑁�X�&oR�/fA4u�4���x���X��@tW�ⅰ�z���n�t˪ga��Kl�f���|k1&�b�E�)&7�(YI��P�k\�)˷
�6�/xcQ�#�2���Q�߂�tOk�ew����V�9<1TV��t�omIE.�Ս����|m��`�R����`� �\�)�]�d�M\�V��gw'�dl�d�Ӎwh�H>��qg�_w�B��yř��v�b��l�����8�N�ec6?3i�y#�$�~E�ߴ��wg�uh�7�2ӽH���S�A�.z`��A �xQKpM�B���T&09������Dnղ�������6����� �UJ�x�_�>-�9�g$���2�6���W��.�$Ad�j��R����x���(I�L|���(��1a���.XI�tHW�H��9c��o0:f���v@ߥIY"s򫷝����3b�"���@�q�c��a�k�h[%�R����a+V=�OHL�PH���-ּ@f�,�Z��K�:�Ia`5����2����Lb$}�Ƕ��jw�P-ދ�"D%NHE��.��|��:�H��*r����BL,�b�:o�~&����.���v���	|��Ϣc����3y5�b��M�%���z��ܷ[j:�J�EF���K��N"hѳ�E�dhB<>��8J�o�nU'X�����Ҡ�t���c�����3PkzMI�3���e!��߮H�eB<����ZQEV#d�	4���QhjmH����S�=�zۋ��dY_�ß8��D��`����9|�K�[��m�<��z�1�W�5�v�Rlo!j�a!^_!��4B�I�=l�>�B�� ���	���Q��m���8Z�9�~�گ�a�«c��.v�	�+��i�D���-�0@[��FcZY&ۃ��gY�4T��Z��|9����$97ux�s�������?3���v�[��ԁ���IJb�ԅ�P�8��~��pI�Z��|"C�����qS�)�i�̩�qj��I���J0|*$��++Wk�A�m�t^�ؿ˵��zڇ`�J]3>P��q��*K�WY��oxY�!��r\�j�}{�x�^l�5,�Q��*g�?�����x"�c�����y�v+Α��#����ZXc��ށrG1ㄨ{���=G^-mF���)E$��{>� �(��8\.�pܘ�W�-x��Ay����U|5Ǩ� �����y���.�)!����J`�&���I�:�TF� �OT󩄡��$��5tE'�9�����jdY�i[�z_i;ۇ~ƃ��=ܰ���5wk8��l�8�O��)�k�+�P�q>�VN��"PǗ
�C/kg���&z>ml�eT�U���M��(�= ���o{�隮HC5J����D��5_�M��|���C��$����7�o�![f��R��pRѢ�F���LBY��G�5z�_Ee�$��i�\	�c�|-� �ڍ���o9!/�7(Ny��C�QB��}и�}rR�Ğ�C��� @�B�2�F؞Nt`ֺ�>�Hv6��Gߕ�vt�|���/O�2{rΪ��]����<��[6�#������h��N0��@����U�������2�S�@�>��΀g��@���&8A �����(���^��(�:h(�"Q��Ɖ�y����!���ǿ�gY]�Ќ��8�6u��N��:#��2�r2ש���Qs��<�ʺ��t�~�Z���=�k�U+�r����&S�_�~u:����ޖ׹�:����b�#�e�8,nh ���p��1��5�w��Np�ټ��!2���{�Dvbw��
�A`�����y@}�p�^W��D��8����M 5,_����CE$�̝���uP}�&W.Ƶ}R%�#���3-e �2w\UsO�-���!��d^v�T25;�c鈑��>����Ʊ��:�`hg)~��C}�������{��?1b�:S<�E_���:������ԕ^F��W��i��ө��a�4wvG��v��k'��h��Q{�u�κ�iZ� ��Zs!/Ҵ��˃�K�Ef2�V�~��C?������Q�O#�?S�v�	A�2��5�}@��Pe�-7�ܤV����!�
D�Q��ni4����V��${�錳�p��f�>���a��~?$c��(�8�?��C��R����|D4/cG���Ω�"ݑGN�_�dpE[ $K5��������=G[��}�.̓��7���j�zWF'��H�!v_a�D"����K��V~F�m
�߽����X�2��Eb�l��!t"����������w%wDE�;DDSs6
m���s2�L?���5�#c�+�yQy� ,��j��B��#����*a��2���u�1v\4�Mc����p8�PO���$�a�$i-��1Q$P	���O� ��NU��Ɔ<T�o;9�Nj��(��q��y���.�gҗs�.��}/�9�5*��F�R>�&�@7�[����X;��C��q�ߥ-�G�������Q?Z;�aI�sq��J_"
��+<�juJG�.=�G�e�dג�m�� ��b��S�X̍� 7gl��"������:8��O[a��;��pbE,M۰���H�)7;Si��w%�Q+���]t�dV��)nM(�mF��B~�qX]ު&6��^	��X������^��t�L/�T�%{Ÿ�7L����R�d�c�V}��`jȭX�4V����GqO������������Z	p�f�5��,K�'i���4<0���C:i�0+0Zu�b|}�~�i5��Ѿ{�
��GwG�a �{J|�B`�(��("7/I�x���<E�_ݙgO������p�Ow�¨p*��-�8�;�d(B@(J�-����55(�P�Ƈ���G����d'�!�`�0&Ջ���6�r�l�<Hb�2��([_�3A� D�eU�`�1����0W�?fg�n������Ĝa�7�W�-A�vi|�]=��݆��(��7z��Q�G���y�v�����fA��9�|ǖ��,���7�'Y��\�DT�G�٥��D�ڷ�v�~u�
�xt�x(����Ѣ���J��V�����k.`�(R��W�G9�ڎ�1DZA�$�}/JM�)��;�x��1J�`�P�.������O��T��$���K����g;�E�g໹��:(��N-�U�(ۅ�Ec�の��ɳH��E9c�(�D�L�@\P(9+XZ�N�v_&�c�]1W���2&����3�	�ƍa�@�{�/T�@ok���{ӟ �ʩAL5����_I-٪����|�󯳫�
=�/i~&�G����B�Nkl�&CT�u�=NS�*����a|̀Aq
)w��6�����;M*õ���a eZc��T�@u�	0D�������M��-��ϟ�O��F��1�OD��.�$�I�C{R�s��s3+&�#�?
$����τU�IW귩�$�֖L�j�H�W���KP�'��έoy,<��x+��.�5/ڤ�)��e�jw�۠~D�����,�J<�Y=��sA��R��}��q�v�a���6���&X��m^���*��ɦ�z�v����̄Yt�>��َ��zj�o,�C��|� X�jN3���{`�0�uC�І���`���?�h�{���;��!ޘ�� R$�Qk�$�BgULf@��D�M�L߄P�|��N��r��K��?�y<����n�._��w�EJm�hز��RH�A�H��K*�@�̈́����빉vE0P�1aS+p^��4j��48b�u��g#��L�#�[|���ɽ��C��-{l�N�m_$�[�ֲ����n]�j�Z�Vc��IT��("M(L��!��>�'¼a��F*��P�b��ޠ.�)-�s��}�G��*r\�'�R�2��N��<_T Ɓz����H��1��d[��{��j&&���3�@�!��
7�NĄ��pT��bA ���Ar�&�����?)l��A��=0�,t*_���d��X��ik>���f�q�M�?:��r��a���BK�/˹���8���u,6O?�t%���knͤI�Vn���UMd�TXFn�K���mp!8��,Z/ŀ������q$MwX�U�%��i�+m�?�^թ�i�	I�\��F��5�+Ε��M�Z�����:�����g��Η��L��+5�"kp--��H��s���l΅
ӥ4���Y��cY	%��j���ro�������$l
��n�}ba�R��bʴ����X]��d=�(�uc>xl�<9_Ty,kTQ!d�{�)��.<�-����Dn�����	y���|�S��cs����ʷ8�6:�˦�E_[k����e��7���#�W�x��2�>�DS�4�7��t����V�8	i�0���o��nbF�Ĭ�<�˟(�9����i/#���o��n��[�ٙ<H1"������t�_/���1t��;�)P?��nӆ>�`��7M�}��)�R�wlJ8]-���6�; G6�E ��`��evd�o�H���@n�}��1�g�r���t���A�z��z�2H<p���0D(	��9*����������ؑ�:o)Y��(���}���/��JS��!l\�o��^	J�\�UGd$'�ŪUS��U���yu�Y	��d�o��耚�4��m�ח��y�Ҕ �R/���wn�r�.��__o�<�61Ty���/�)~G��ki�+Gg87�b�;V��#�$��xn[���|_���`ԭ��u���(�DC�MFlAp�^$����P��c��߳19IY�4:���w��[K�'	�����)�V y!l;�l�s#��Z�;�碣�����&���K���A�ok�𡋰��e,��..0n��,zAoiCO[m�Ő�zclY��w�|Վ6�H�4�T�p�2���4���s3��<J�T,5��8�1%o�%H�ʃd͖\�YKc~(�����y`��T%��B��0L�#�U��;D�I�9ԀWՑ�VYm�z��N:e�Cw�`�
�)�.���ߌ֬��18>x��Δ����6mY�a4�Iw?��ةїe]u	�o����ۃ�ؔ��9g��j��³K�����B�lMDP]/�]�?~�*�d2"�ն���4he�>%.���W���ƚ�U����<>�!B����M���xt4p#h��LJ�5��?�/�T_���7~��1�q^�^u+�l��9��I��^*_6��,�ж���?�}y��I�i��ˉ�ɟ�R!��x�K���-��"�Z�,͔����r��h#�~lb�<`���֕^-L�xkW�%�b  T�IN�1�
�r�L���Pn�1]�W�'�2w��!h/�H��8�Po�5Pk	�P�N��d��L}f��3EV�#JIӍQkpݡJH+�Pb͇n�B���:�޵7&�zY�V�?��A����Ʒ��wd�00�������C�4t����Bޝ5dorm�b�嚐X��bX,4iXQ�Y�*�k`���#k�`��lt�:��L4Di�W/���[���γ�A���H:��b
���A���NX;���Kl�ĕu'�.�?�Q�2��C�p��%c*'*~��^���<f�P)"SC�[l��:�7S�[ӑ���t��?�h
�1�P[�]�]�B��qȒnGz
ݲ��ǂ�0��+c��ۆ�ܧJ����c��]�|d��oڢ���i&�����A��u�!)RK+���ǡ�<.:O2h�h�W,�(�X�j���&����՛��<Q��'�$@��R\x��qH�%<�Ԡ�.B�1�_"U�Y��%����S���d� �g��rx�|�-�:3�eVI5jw�XR����t:9J�ߎ(��kW>�q�C��2,�6�&��U�����X�/g��=H�WYS#�!/{��BXlxVHYEB    4f62     b50F���PU���t90	j�2���YV��DmvZ�/�v�`�QG�*���l)��p��-�!���Yl�J�
΅q[�3 ���[�ʓH�{�bg��f�TG�� ^::Bg��gN��a{[�|뺅�B�Vu�h��C���
�,
Wv@��Ra)�\]-�_O۩�a��W�~�F$�tU��a�����E CgJ/����L:���3�Xi�T�9��"M��<0�N�P�.���%�4	��I�,�|���f��+ٱXeF�8��Tؑ��LF?ub�H�^}%g�ͻ޼��$�a ;Vl�G-+����e@�����G�f^��t3����r��[�=�hP�1��������i*��~1���2������o'�I�� �U$<^�4�-�ϳ���$߰3��x(�5�Qw����m{�;R�B�i�+��T��y��H'�s��<��<��y5lq�v�9�DN��4�[��[��v�t,Э�.oO�
n�I�4,_�ӣ�I2��:���6�vrۭ��v���S�ӨG3��}۔Q���֟������q+}�G���c�)�Q�5��Iڀ�4Qs�L����O�܎BuT6��_n�dqj�N��;M�_���k���hP�?����*��'�p5�^Bb�*�c����B�n����I�V�R!O�A�'2�C�"��[+Pf��h��ff�ӊ~�J����<�ěu6�c=)���e>�A����2�������O1��!�@6��W�vG���f�5m���6P�L���������I�P���V$F�@�K�5A��Cl���"��w�{�_�Cz}^R�Sd���FN��Uq�,A����{�6����K3�����r��<_,02K+ǸߞRK��1��L��җ�]�ВI�V��}�) P$��ָ�KG���x��n�� X R�ȳ��謦iXPF���h*m�B�o�|Z̉Lռ�''��%fi����]Q��x�Yx�1-�*Ja*�6�y���^ha�8��4x�G+j�\]����{͉=�2���F9�*vX'�A��}؎ƲG�N�5�e���ک�FH?����i3�Lgg�M��)ŬƬ�D`/�qg\�5Ф����\p�(o�s�i�"�z��oĪ��;5�=�f���,���#�N��/	�f:��n9��U���V/m^i�yO���&�<M��k�2��/�=
�w� �mcٸ/��i�
K���*EM�.�B��lj�ֺη�,��՗O@NK�,�J@U ���︡Do��Q�}U�.�}Т^D�9,�kZ4cuN�L�Y���31/�-C�
�Z���N����Q���宀%��'Kū���=� Վ�KǗ�(3V7���j�8�{Ι��[t7������+�GXœ�f���;��B�.uh�i��b6S�oיU0���b�p�0,� ��1��}Q���q�b�vQ�����o)Hp/�O����H��Є�&���(�{r����G+Ia�+����/�jMlE�շ�gc9��A[]Ia��+�'�e6/VĜ�b��Ŋ�j���F�?8T���G�.�~)U�f,�k�2Z'�
������o��_��.]�s.VpRL;\�g�b�Cɽ�A'N������l�A���ĸ��(#W��۲M�9hrB�E��2�T�I1���̿z�u���U6���;|O���v�+���0���!t�Ｂ���T�!P���qcgĹ����w'�ԡӇ���j�!������0��̈́X]b�p~ky��$����%M�<�8�a&��>� ����M!�B8zA�O��З�De�e���B2x��-�M�S��h� �+�3������3<�����hߵP����!Xc�P�A��z*�\N?��{E� �;�R�[��ۂ��*Y����H  �I�� F��\���X�� �����b\�p������=�w� ��;Cja�Z�ZgDv�F%�z^��_i������h	C�g�ja���'�����yCG<�-�S$�~$�J���n�%b�J!0G��OB~y��Ƭ%��Ҧ��}D��:F�S���d�Q#���'�ƛ�ŝ4&9F)D�ȂX@e�|��7G�spw�+��J�֭+ͩUy��:x�⥉3�A�*a���b�֨�t�I��
��yV��YK�N�������I�vQ���]&��h?1�⬌�Á��͸���R�Z.�4�bjL����|�**s/�jB��cNGn��hS���VgQ(�Y�AV�����qй5J#c'R������2�7[���G_��a]5.#���l;��6g�ؠ�!:A���c�mV�9�&>��K�*��A>�J;��3�cҸ��.���$k�}��"|�[9��歎ct�]X|z��3uU����&%iDD����Y�R�Q�%�aHNp��κ������2�w<j4����wq�Ae��N�+�H�ew�����v��ta���3u����>b\�ә���d�㽵�ŲR�}�({+%����0�j�H���ߘ?��}~��RCAƮ7!��@Z pOB�it�1ϰB�yu[���р(I;�����{u,`�,�-a�Yo� }J��1��tk!{�(`��F����[� i�k�u���}k��k�*F,|[o�_� ��

8�#�m�.����4F��-K-�q�	�7t!}��wEx�5[�\h������Tu�]��@�̯�w(e�mz<B�d��j��}nSS3[�LhF�Y�H�嶉'Զ Z�xr�/P��O�C��W <XL*#�3�@����K��3:�T��VͲe�K�LD�[�B���]�a���@�4J+���:��βW��#�e\�F