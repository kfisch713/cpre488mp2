XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�ci�%c���'o}��_}�7˫���1q�K���,��@�݇q	��q��-��i��^m���F�S�H�|׃(C��������)�N�f�m���h"酪�i	����wRY#���f(0e� �٤��Ӑޱ
�����Gݢ2���]xV�(dNzW��V�?��n��i!����\|v���D�Ds�@x�`XK[(�k�38�OW��w�i��^u,���,�����c?��P�
*!pFB�p�L�	��9��+z�.�-�X䥌�U�)�Ο��rE w��(�P��6�q������F^�ZĠS�"��"]��O����E��/��P��)�0�4L�~=��q������L��Ș�� �Ş�ۀ.A$0�e��mF#L����+�����x��]���hb)w�D�
M�z�E��5���`r�������L
�-����Y����.hT`�� �Vb�W�8�����nl�lj�K�c'qk�N~2���9J���n���u�˃�1I���V0kg��n����R��K�U�~~~�4N�����ӕ��Kų���6;�o���zJ�#�ά&����T��bdԻ�ho�
IR^�9/��
Z|_+����d�[���'�	x�Yq�(������ሦA�|k��	�职�7����͊gi .��G;}5�K	�7�3�tlX��|�Om7�A�������&P�SOb���O9��ȋ�y�@��X�R�㧹�>X�7NH�7I�XlxVHYEB    3fdc    1160O�j���tt����/@�{3]D�e����WU�r�į
�V؋=ȝ�(����
���w�'����3���W��;�9���O��u��KU^�^�=�ОP��� ��8|���H�T�'�LX�*c��!tf�h����v�o�� nβ��	h�SX ��sg��2s4�k��@_��/Ae@qU�)U8��-Э�������t����/������cວ�p�xޓ�k����e|Ӆ�1���F�i��?F�K������>���]��T9c��5����(�gl%h9P�	op��Y~�@d�p�6W���2�Tc�j�R=p��/���Q�LT;� �AE�[_���|ݳD;��c:Xt$�Uc���	�L8��m��d�\���`5��\_B�����9�쓟����0�֚�gyA����J>E�Y�K��*꺉��7��cC�1_����2B�*{CYL{��ɨ�Z�l��n��+���S��sb]�7��,\� �"��Kb٩��x,�'��(>g.�4K��{%*e��7�ׅ��	���غ5�*���Ô �~^%��4H�)a��hhw��c�	�9�����z\��B1i�BhBa�>�����p��G�+�쐸uNx������'̫���И:k�Y�o�8�VT�Q���*��ї�#�%H _�zA�D�	]>�N����h�T9GH��۫w����p��C��Z��S:8�`�������K���TB�q�s����J��-��yByIb��7��3_r��
�<�̏-H��Q��5W%�c�<�{^,�佰���[:ધCP�l�H��:���å�@�mK!�n=�y.���s��}���fy\���!�3��,I�J�1��t�F`̬
j-\�xZe�e���(e�{0��b�Yɡ4���.瓒q��= ���L7y�9�j-���v�=s���'��>��i�k��/���t���A�-S��"�~�3 ��6��7m��됧$�?��rQ���T�U�u��j���`���w�Ӫ*�;I�?�]����q��?�H�d0'�Unh��%/�+��ѶZ�k��9R��Ϻ���yv��nY��5�[_����z^�ו�U�L�'Q�1�!a5���Ds�������g#����6vD���H�Ō����7�e죱�ќ|�͎[;/���xͤ�kяD�O%�W�Œu�^��Dem������.z��H��̌�VՋ l�Zz;H4�n"4�$eӫ�ěL��bfsS��q��@(�������Z!���%��%Q
�$E���P�QHSR��!���RJ�+;tY.�g��N�*&���3=	kj2�����=��7=�&��}����1�W�:��P���Xuu�L�D�k�ߦ)'Co��!pJ��#�ab1	
7
�"��\Yѽ)Y�b~K�ڠ�>�5�4�0͑�v�gI=���[���,�Ai�1����I
,ן±��]~�$6��+!�" �Q5nQA1-+#�#k��P���]CkI+"��$�F�G���ߠ��M��8n��K)��Y��A�*-���*i�1XB��.8/�뷧�W�Ap���H�s�C_��(�F��t��&��!nfA*W�[�ʸ���u��n�LO�s��?[MΠ{�{sD�H��w����#sj�ȆJ����N�[�vH6���m@:+=�L>�@�W[<�����BV��l{rC2[���^���) 9�fJ�j��]�˒쀤��u��w�*\w~#(z4��-K�}p����Ze�R�Y�$ڎ�~�*��$i��vs$V*C"P��5��_����w<�	���+��܆��kk)g�bk_E\А��0�#ɂ^��!� `�_��Sr�'%�a�A��@�3>����a^G-���"o4ٍV�o�Dё�y�I<-8���
������\�o��^#YFg[�f~����gX�_)�O}�&W??��/D�&�A��-xfd��i-ȓ��e�ˈ�W�W|�_R��w7�1y=��f��P9%8�����pw�Nu��4�ᇧ�>7 �uq+,����؎��uX>ǒ�m���r����$,�e�C4�Kk�uN�7�ƍ��i_q:p�$c��E?�Vv�@���~�"�/�ы�s����$�\���U�=�����-��
��pR�i4\���ȏ8���q=$hب]� ߃_(q�pێjg�#�w�f_R�B�:?A�%�}����8�bH
枸��$ʣS�g\^瑄d�E%�8�r�k�e#�Y
�ā�~�c��1��46�g7��zG�}�V�~ЩsL�����H��QF6H枳(����b��B���\�,H�b���sJF�̫�1�
��x�i^{h�Jw�h�5@�-HY�B ��l�6��*��刟��?,*yH`xb��7��&:*+!� q�Ks��F�[���9n!4y#�!r��jj��28�-��6$nlE���I))�����]��z�ݷvo�
s�7.�dF%��^}�),���!J4��<[%B7���0ڊk܃.����a����!!�E´EI��a�S��^���=]u�C�e��+?����USe�t��0�"�G�� ������<@b��Jڍi�K"�u � 9��"�Ο�2v)l��U��|���xu�__A���c|��XI�z&̀���:�^AV�ȝ�D�ORכ�{��1"��3���И�űhRςԪ��v�ofQs�0cܲMp�Nڍ<쒦6 &�2T1�6�i?=x�M:�@��hEߪ@f�H_�g��ҝ�~�׾�>��9eܤ�+�p?��Z�.$��A`<]'I�:�t� �i_R��ͺ�(^So׭�3W)����v�(�};���%�������BtT�H%5���^���4��FR�j��i�ܗd+�!ZD��5C��RG�+Ͳ-%q�O�]�c%}tYW��/��L��i�J����b�j{aքb������$4N���Yu�b+L� ʷ�l4�9ʕ���xN4�e.���l�.�ScO�^���vG��qI�ڔb�����^�%-2T�trÁ�ķ��Y+�.vm�y�b�����|�vyL�I��D�8��"�6�a[ �>C�O-L#e�>�%uO2��x���Ro�"T�'��jW���л��޴�VQ �r>�.:�X�������yV��)s��[ �"!N�R�Xo%�,�,_���"�� Z��@�ywP����t}WH)ڞ�p��i�#��N٢E�%N�_F8Ѹ�?���܂o����:aMhH&�D�����FK�$��y5+Ȇ+�!%R}�&�ƝV���Kycj-� ��+�y��*濐$�K�������n�VB.4ZU�w̓�h{����z�2]c��/[����t� 1���#�^���}��I/fHd����n�t��Xcg�銏rOx��z;[S��j��wK�T��|ncѲ�(���x�<* �^�..F���^�u�������tG|��7y+s�9j���l� rݳ�:��N5Y�׭���%O�+�)��쀆�v�߾��IR��jI�������VG�30�e �N&�@	�W#�΅�8�$��D1�IR�s����e�m-ϗ�ڋ����bʙ���*+�Cg�R�o��L�]e��¡�[l��T�u��(�� `� �n��$��gBP&�=��B	�Fv�ཥ͈T�fr]�GdE��(��ޮL����s�Z�ݦ���4��)�(J='�nks�Jqe:���?u�����p�ѩ�K]ᄝ��n ����U���ܒ$��	:�B$D��1���s>ӷɉ,aM��_�R�4�.�cW����^R�c��=��*Ik i�5�����郦�,K;��S����J}ekGJO��@nL/��������Ҁ#��w��6v,5�sAJO k`�H�󉽘V���V�M��i2��@�Y��� 	]6���]���?M_5�K�������,�u�|����.��"��<�66[�P\��M)��3��Q�f�2��R0�:�e�o��ptF�#S��m��ʇE�����7�����!��h�*߈�@=iM��+�	ggi�@��;т�z�µ"Y|�h�m۔�w�ŷ����
��?M�9�JW>���Af�BT1I2�����'[eJ�[�.��=�Aְ���(W���/"�V�qV��zj28���M���j����S�X��t�Vʦ���nX�`�_o�e��kɟs��{��ڒ�2�Gv�O�Pv��!�8�@;����wY[Ǭ��r�a��4 �5�U��rL��m ��^�y�L4	��!���@!� W�6���ʴ�U�~_��@8��T94h�y��M�m�����z�s��m�o͸:>�t��Q+����=ر��}M�'`I���#A1