XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B�9�x�Q��n��|�
mC��ݵ�C��}���'�in�,Br-1�K���;W�~Z����à�g?�(�*x_ㆶJd}�#��� ����I�d�^�CDr��3���g]�᪭J�ϰ��cV��k!��%N�x���%�=�nθw��,x��  �؂���>5�q�ی��+up�����|;��*u+���q<΋�5=F���}R�_bS�
�e�i���/<���ϚDkZ�]@��M�p�8�c�P�)h�1�70Ui����c�G�	;LXN�X�.�%5�beM�������L���M��-���L�	Md�"b�&���[��T�f-B��K]��'e��xAc�3/�\����4%��>�6�ŀ� �a�׮9�2!B�*o\Z9���Y|J�ό(�L��S��I���	��F���:|�7��nsy�и�������2ƹ��R�M�&�Ǵ��I�\��/t�,/�2�
pm����/qȿ�E"���e�T�0&��A&�۱~d�z����7��A� �X�U0G.�.�gX���1�rV=�T ��;����n���f@������/�{Gi����Df�<�}��錏�i2�ϓ���W�j2��YI�[ڈ�ɖ��W�����s��j�ߴ��D��|bʣ��p����)ݦ! �a/�۫X�&�����+L�Z7v���\��G0g��� =x��0�����I�$�V��3�3�59����%l0�R�+��MWfB�XlxVHYEB    7265    1660�;RR��R�SڃI���H:���	by�w7��ܣ���F���f��/]J)��w��ؼ-ga��z�3���A��]��K�z5
�Rg��'����!�I�8E f�B�4�M��h��3�{�_��9NX�o�G�1BZV�uM� ��3�wg�*MB@̴G��ճ}n���Y����e�� �e��*�8��Ջ��4q2�Xe�dC.�K����+in���u��PH�Qz=p�aڷzp�����oN��*I+��P�C�q�h�1Q/3�0r�����8 3��!U������<��DU��8�������S�������x�sT�������<��:�.,��Z�'�X��?uF��z>8�����/�8�љ8Wy�Y��:�Ty�7w�}��aAR�������z/�f�ʸVCW��/w��: �r} J��~�'ۏ�y[3�T����@ɒ�2Oy��mg��ZP�*3�.8x+��dw����i$���S8�*͒�Ϯ��'�#���lb
�w0B�$`U�P�u���ƫZ�:$I�Q���%ll�#�d_�v	ᰚkUm`/GLS����%I�p,+�A�$����5����@�����"9�?A<v��j*��~^������r��p!|Ɩʿ�w�X�����c)�i��@Ӕ7���	u�'���'��=�o�Ri�� ����Ʃ^2k��J�e.p�N�+/�4��ʫn�	J���L"�ya�}9��u�3v�W�^T��N��[ˠ+�V�ㅕ�*8��	����3�[�Ԝ�����B���Ά�.�
��|dڐ_���ZT��v�O6)�#rG����o6"��ϰ}�3v�=���3r�r�j��ty��[���-Y������M�م��N�y�i�4�����ٳ6�X/�bd֮k
��8"w�U�P�-���A������̻z�� ���3��`�E5�W~��!
P���
�D�Ga*geΥHC-8�E��6!�1��1)J$z��c@U ��S�˪�g�Ӵ��w�2�>�&M}�� Ҋ/� �Rp�)a��6eH�N������!z���^`�_�n(dZ��ސ����e�Dg`ȼ(g�B����s}�u�o�y-�p,3.�!����ɂu���I��ע��@�8Y�V��u���%��Y��@�����G��A�Yr��<.1��c�:@�:7���.�{V�g��"��:�5NT��xHCO��!me���^�	8�(Q��h!�F|�UK�+�����%SU�/�QQ�سGY�����;r����=Æ1Pa&�ZЇ���D�,����n�`q��)'g�� �X�!���+��Uao��?�����g���1h�t�f~̆�X0I����l�Ǘ�~��������0���F�����8�&�%�q1ɭ;Gѯ�
R���&�~C7r��uR��$��P�N��N��V��ܰ���j��v2�h�v`��g��I�|C��OSԂa���%�a�I����gx��䬧������j���K�ҩNk��u�jz�ǇL��W�}0>ZD���])h;62\#�[�����_��3Fj��������%�A!p\��7�c(=�t�,%��%x�5	���~��|����
A��|��O',8i��p�cm����}�_�hw�!�C��l���Յ-��t�U�Uh�t&�篊�}�?p��� �K82�KZF�P��R�.M�|~)k���n5%С�T�>?���A�f<�~5F7�s��)����,OY��l�G#!�'��11{���e��x�p{��W{h�'���g0��}�x�u;NxF
�\�-��>�#o�ݳ@'?�jC��?ٻ���+��~p=뗭R��h�8�;�.��8�O��%Z��2,`4(,�@��X�! ��t]^U-A3U���}���+)�BP	�K�b���g�)Ȩ$�E�s/��?h�I�J2��3��@WE�h���KZO�@B�Mh�7�z�[Bɠ�I:��l��\B���r'$d�%Ӄz����0���y�E����:g.�Q��m��LkCz��P��k��m���S������kd�����V�����������@����:� ȕ����4��D�Snz���d��ߞ�S�h�x(%��)���M�ϫ�XV&�ZD��*�$31����N�}o�Bִz� �p`pjmS�xς7I�����U0����p�qx�,�0�w�>�N<�7�p��zU*�McvD`F���T/c�Y��=������lpg��=�Ck��yo�-sKy�V�|�O���	�+�:�����u�
�9�pEU���hP�kҭƷs�dbi��b�c�I�3ڟ��nu�p9X��Ɨ:��`%I�L��Wt<}Of<�䵳Q�|Z�eg��������U;�\Z\,��*����#���o՝oS�s>�/�C,�'\��8it*�N�p��صZ�M�@X0�J�a��W� {K�>壉�*�.{�b���o��0<~�\��Wų� Gϒ���У�@=o�[�] &+���#�3���m��B�J�R��k��;w�ٶa��Ҁ���h�	�61�Lh��j��� �<�$9JtP,��.+鯎D�f�q��eV|��N�9]U���p���9�S��C��3�/��'�}/7ұ.ꢥyQH�ev־qv箝�.���oK\>���b%W��z6�Y�ꈑ+�s/��B�W�SN\�iR���,�ց¸C�H����u(�Lrꂉ�࿆C!��>?�R���J��^�}{�,8� mJh�������Q'B� ���p���ii�>]y�[��	�T�x��g�uD��Y9"��������*C�گ����Fi�`��Q�K���a�T� �Up,��p?�[����e��y��A-��QA;�>��w����Z�GؔR�@u���u�:*�`{��`�ʉ�N�=�xM�N�`50�(�����+xbo���c�x [_�~�$>���jA�gU�k���0������/�'�)n{���r�KZ2��'=\��y�A������_d�Y,�ƛE�܁�m,!��6��bfS�w6���k_ �_��a������KP��AA	 �4@/X�[N7�p�>/΢D?SK�8������ &���� �72L������3HZ۞�9��;��E�����������oR�&���ʳ��N��N�S�۴^	��菂u<*���0�����^�6�ۤ,�P�BF�C�З��FzrS(� ܕ��|�@U1(���,*��>7�}�d黰U�����'�;����wX�Y3����/���Gu>�����q}���ڣ���h+��|CT�#�O�E!o�~qޕ[.�-��O�_�)q���ǡ0�T[Z^���),�G�LTd)��x&�y�;��cW; J �\!�� ��g@�RY۲CE���p
ԪM�	��#kX��lε
��P�/��t�u�*�/�X"�$���l�����<�](�b@�/~d
��Ms����<id����?������鈑�tl�蕤�7p�?5����"��P���������dR`!K���ߡT3s�Dwv�vSOx����"�4�E��>�q���81lϸ�k2yy;��)W�_;3a�˲����8�z[�I����4�"�\GE8G����2jv�OVƠ{>MOL�H)���w)��ʒ�ռ+,!�[Q���W�R�դ�n�pf��UE�a�����q�"[x3`��2.�uZӵ�����8�;��#;)���7���vZȬ{pGiz�@kղp�gK�,o���g6Z���LI�v�,ay��H�V�=3��=�@�}�5w�
 U���Y8�>q�#.��(f/��[YPv�t{��I�ؽ a�O�W�8e�4���/V��=��o���;�hĻkރ����fB�F�Ԗ�țc��Piv5�xtE(+�����G�`*LVᛍ�����ʡ�y�^�
�.�4]U+��6]�E�B<FٙTI���&g�;F�!���LH����2�i�7��1�ϱe�V:��@:�3.8`~;�>L8K\�V���ů;�M����睐`����p$#�)E���楁��c9��~1@�=�0�N+p��t|5�	�_����%����(c2�7M�O���9Ɲ:h�.'1��
?�g�����Pxt�0�����)�*�(u[i�;9@Y��j>uX�J(����В�l�ҥ����0<�+�*h�jM�N�e�,TB����.|�k���vr�9-�UG5�l��M��],t�,������ߧ�2������˙|�4��!���l����+�j�fZ��A+�&-����3���n��޽X�w2��<P~�Q�$�O�GK��ɪʥ[���vr 5�Ѧ��q����t�8�-÷v=V>�"-�ZӓoX��y��*%[#2�Ӱ|�a5�:��4�xo nMSī7�9
r/�I��^(�e���K�2tֿ��D3�6DFj��A�N__�%���#.��"oZ ���M�D���Px��hX���1��*��}�&b���V^�Yv��OB�'Z�cQ4�<_���S����b��r��C�{]�@�jѸHM�N#JJ�B��&6��+��%�)���G�8H�.��q��)�~W�DcAPS���סT�8�/�9��<�� �t�
�!��r��@���	ѹE.�;��"����<�Ɂw&���T��Uq����S'I	o�A��QdM�` (�Ǚ��z�(�+}���Y@I��g��Á~�
iQ+�%��K ���s���b��z�g�e�Ko�$�pɾ���m��塗�ֵ(On��H�P�{=$t�� 7��ǘ$�1iLZ�B�!j`��JG@�Jt���`��cƂ6*����6���6](�x;19�+$�_�2r��J�����Q�T�b��L���$y�)[<���Mʒ�U;}���(�xʼ�RW[��0�G)�̾
�)��F����\$.j:Z�� �߻���[ppO���UJ�ϴ����oe�k� 	奛xѴd�n��.S�pY��Z�Vl�?Q���M�`����0g%w��bX�����:ț3�q���tB{��Ik�&�Řs�8d�{B?�r�����@�� �o<I���g!�lL1B����K\7 �=c<	sg�Be���dQZ8�
Α�:t��hB�D�P`~e	O|�����PTG�C�L���2e��?E[a��S���t�W��u�����j����>��8��{3Ջ���)�+=�Y����^���y��B��B�oE��x�Q1�f�-��.~��䟎�a�JvY`�%�o�;��H�jl�H��Y�R�t+;�Ӳ�0=3|:&���N����Y�/z�/����Ȝ�����*�E���Φ�=f<r���R+@}�W���$�+cJU���~������Q1�����Y�?��{��Y^6G�%&2��?).k�͝u]y�;Z��R��ە	�%�d�M��P@#N@�FO�L��z�6�;�T��qK &�=��p��fd[9B �tbﮣh𛸙����H��KF�Ҭ�^�*<(�n�ͤÁ9e(��'���^%I�,`/eՆ����'o�O5|
lĳ��l�