XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��qk����WJj-7�����i	$�`� ��Ҕ�Uh���!������������襪/|��'�3��=��,(��	D͹d��j&�D�[����;E���M�D)̄����9�,��%6�3��8�.p��v����|%Si��FĈ�/vq����5G�&��M����X��*�����,4h�!L,-�|����m'����Q�^3FK�dy�ҿ�U�R�mw���p�� �4�Ă=��A�n��I�Q�mw�?�0��jMCy����L2����9
��a9A��:���˔V�3�27������	�Lf\�`��M��W�s���M� ���`=�+���Ny*[���:[�Z�l�Ix��b�L�'˼ZǀRV	x�nM��F�m���ˏ��	����2˱��B�of�Թ��|ȶ���������3$��YT�SL�LH�>�a����L(4�8�������(�<��+�c~��ԕ�/�ɠ����D��h�i>ϊVV�A{(��0C�������R�	����PK�U�b��ZH-�Ѕ�a�
ۉ��*$ ���B+�� ���s@�P�sI[�����̋��Nm_���9C�˸B��7:4��&�Kі�|�r*�CP�v��>\�F��d��Pl)��T�>�gKUzm��@�GO��͕���-�����1`��G�����go��]R��XT.toq���^���9�q��T��)�M1t)�̲�ށ�_�[�5P��`LXlxVHYEB    5224    1740fʠ�RU�CNa��M�X�{8���],X��5&Հ��(�4h��be��VOt�Z'u�k�%���/��Q��	=��%�e>�L)��
����a��m�Q/�0�.7`3� ��|��{� `��b��s�w��~�+��G'yƘX?��C&A�v�ڿeO�6��韥�����r�y���Y!R�Hy�pj�x�����p�&�<k.�� �$#�B	�>�K�nN4-''�h�H~�ێ���q��6�v���� �ʡ���s�&+l�(�O%�Q��Ԧ0uʇ5�'�Ѕ��H2��%F[>���̣C������&���;:��|n8��um��Q����2$�V?j>��w�FR-E�����4��_nH�8�w&�Ap�9�
�ļ4t��q� ��yX,����(�3�&��K3����^5�6=��Jgh�Pi��2���Ě��9֦ ���9���/E�[x׋�7�~�hA�D,^�*�oY�a�s���e�UA}߷�1=ڑAgDƔ?�X.p3,Xˌ�,r|�䌻l�y� `/����%3z��wV��Ir�Ģ��AM��oA�4}$V?����J�(T�u����1<�Q�����*|W�����?I��i;�F�X��p@j�NF��ve�Xi�������j��q�'�>m��?�;F��Bfc;ط�o��d�������ԓ�R����LY��~l�X�:��Cg�Cy��rR��E�#�&՟r̘�'R�ؘX`n���� q�#��G�Ux�����E�m���p�jm���Lu�OÜ"��(�e�1n� �g-䩄�h���P�`JwL���@�(F�T���N��W�+�����5^9b/Ңl���c�7�+yƺl$���d��U�K:��-����T�@~�Bc�m@'C*~L�b�(��Z�u�
�����'1�Ll2��W⭨��zĝ7��W�}��Rĩ��nh���&�D�9a��u �!�$��oJ��´fT�� ʌ���&v������1M]�~�;��̦��I+�ڂ���Z6KW�&�~9�p�ޤ��TY�D��	Y�涗�ԯ�d)���jI>X%���j�W��^��Ҋ����2�^������ځ�.����o��{�Da�Ǐ6V��-��;�3�-�RL�s��9�	�Ku�����7�g��e",��A������H/���$6C�E!���	��u�:��׋���<�6���hd������;Z'�����:կy�#�N��s��7�+����yV�,�Rd�1S�����}�1z���>v�#h����d�0*2x+.L0�����C5.�?U�
B(�����6S���~�'I
�%^*�h���D��}%�Z2���ͬu�$�픶�"�4����0\'�uu��h���]�f��Y�*��0w��Y̑s������A�(�b�q���[t��v-OYZ��h����'����5����
��c#�_�3@�����̕��'	Ϭ?��͠�`�����7�"�U�54ֳ��}�k���3f��c�r��S�5�����k\1���W~��PfxT��C�_�@(�Y��f%P0W�!���EtcZD4cc�����y1x2g��A� �p �\�0�-�Q���fEl�WqA
E�G_v� ��1Fd���t��R�3Pz,�������Ɇ�,7�h�\���ѩP��v��T�R��FcGX�v+�c*�q�71�y1�8g#y�T��
�?��#�I�T�KL���@�1�\�i���2���l���C�ʼ���q:�O���Ac����f 4'����S�D��:}�Zb�%��Y��mR���n�ew� STW|�`�R�{f��W��?^E���7�Cw��Ay�k�ꩩ��P�5��nm.�H�D%?{1oq�ØN�)G�~;�Q��qE+L� �I���>WIh�����qb��S�i�����/��Uz�����M���ͯ������]~�8���Ы�q5���!~V�$V�L���AG��w^�2]O�����(��I���������b�z�( ����9U�V#�b��$�fW%� ���rk���@���[�@\��z��QK+.��8;>�[�n�i%�g YtutI�m�v��s
�9��*T�$��vxk��.��_�RQ�{B#��\�����O�? W�m�{K����O$t�R�8J�7c�l�1�d�I�Җ�O?���2E]��n�p/7�q0N+�6r���`�~c�Ļ�Ai�>�=�$�pw3�j7�8�Y�ߝb}��E�/�w��E�d���\St��V���c��t���4�!�z�m_`��b6�>�ãC��sQ���fd�U��g�sў �*8@둹�y�lG��61���*�8ċU-���^(W~��!�i�_�n`�; i0�=0�)�#dE���D�vy��8�u��`f�&)H���<��O��2��;�hQ�0as�����=�����ɕ���J[w�Iw���h�y���lk
|%yB�G�,�B,���)���>&���W{�����<Vق��iLP�T�k�k�/nē�2ӕ�\��,gK�a�R����r稰�mAF���:���g,�F�,6.�d�f�N,���6�#�Y���^���*~���
��L]g�5�x�+-�WW;�Z��i����	��=�n��G�2�D�F�C��ݥXoOG��C?���+����yq^�U���9j��M��%�U!���[�ƕ�� �Nz��qK�(�@��H�:l�J�%�o������ <x���x=.��]�ّ%�wqR,��R�M&%p{c�<�6c������`Ga�h�m~R+��z}y��~Z���/��=�oӘ�L�A�n����CP$'�#ھ;�$�
������(��s�W֝���բ-���Cp(�^��3F��S�A���S&��6yI�-9�^ף��|�W[;~t�#�l��K����=[ǳ� ��i/1�5�M�b�Q�ꤋjH�3�
qm��?���:�~ﴼ4�n�*ߖl����?�BC�������5�td���	����z�qGf�������J}�)����u��'FB�p>�G #1�4
ˆ�ψ	_�����6/^KsE�c�k�x�B~���\��#�.L��o�U�q�n�`�1 a@@����m���m����m�L�W�,ѫ6��QAM&)�Y_���dw�����
¤����s��k'f��04�L����/���1��A�����G;�>��Nbo�F�.e�����!2┏����q̯��+p�;�f�;���yo���u���f%�v�U-
�ϲc��f���i+F̉a��Z#���'��9�Y�A@"`�q���M��v���QD��������"U�)#��'g�;��nd���'�KŮPXSqM��Āl;�H�YT^3�[��6Q['%JGn�B;(�T��r	F&��$�t��z�|@�`���xlE���.����M��|�Vx֑[ҩ�̯�`����v(-�g���������! �&F,EamKU���b�}ճ��򊲁.H��=cW�7 ^��� �������PB�&a�k��hE p!�.���G�nJ��=)J�a��I�������(����/*Gj ����"��Ц|
�2��#ldT)��Ե�ԠJkh����6IR@R[���*��	�IZiI�w2󳧤�� '�eǔ���kl���W1�uF�����
ٜo
l�N3�W������"ݕ��<7�L=D�]G@��f
s����������:1[�.��]����2���!d��Pc2A�4��'N�V���:��Q��l�s[{k���2�u�?���	��~��'�@�w=s֠ʊ>$��Z֓p>^�(x��*pn�%p�X�.Z���y�HJw�s�X"t��&VG���UcS2\�վ_��ux����U U+.#���v�Bc;�iĸ��0gb[|O�+��h���ÁD�X9J�r�C��ȫ���y�C|RNNvIwc�쯇��a�<Q��s�k�@U�q�� ��*@�_���Q%mc|x�G�~_��A8s{���q��r4�7�LS$b��{D�y�4���"��v��u����8_�R��c3��:K��y2i��*A�E,�8��A�̀����Z��%Bse�~�c4� {F�UM��M8�4�QM�⧲b��NZ)یvo��&f(�������K�}Rp��[��2��g�C��ҥ�m{K0�;p�ތ7�i����=�H]W߄�n�v���~�����g_֞L��<o���u�����*�m:*h��NF��)�0nmĞFO�{1e�a����C �a�IHA⽘A3��
P�=3 ��B@�i�I�j�)��K'��� Q�aL�ʹQ��e�5B����7t�����:U���M��L���R�Y���zU7����6�z�%���������W�}]È�36�-$�x������α�+�=��9�����]��"
��>�f8��K��ꃔ�B3�>�ݴ��R罼��yw\$!���Z�93��x���xw��0����N����U�����(./!3R�Q��qH<�OԃF׭_;%���kY5���KЦgJ��vm�V� d����#1k�^�V!�K�K��f7�C��l$9_�{@�͕�S���n.d"$�צevR����pQGʧ��;�z�a�M]a��y:ca����>�ߡ8�HivU�z��H��M9��+�tZ|FJ�oS
z� ��:(y���+���䓅�kئ�5����a���/8��ݤSs�TmIg�N4w]��xʦt�n�cc�U��f�T��:�(�ҧ���:~�*��H?!x�ajH�թJ�L��*#�D����),vcr�o�{��P���Wx. ��=XϾ�?Y��=>��܄42͞�b���,N�4qSL�F�Dq&?0W;%���?wr;W���Ǡ�	b��GB=�3��r[��;�m��'Ջ+���b����I� #F�){jV�X=EN��x�C�[�A>s[%G���Tz���L�i���&��#�4O:�?�+�t��b�\�0 >�˨���ʼ�|�M������	��&۽�X�nŀ������)Θ�O�ML�FN�5$L�t]�]�z��{��a��O��S�\�#w�2�K�E���Z�7��5�r~J�"�T�');'�Ӕ�%��G7Z�+�.�������2I��Mmz���&Q�垊��rޕ��ʛb�v+����[��&c��L������	W*'���$$��M D�v��d�q�(��R�0Zu������=�X���em�x���2Q��X�Y���m�E�,�]�z]o��?�!�F7������CE�P�����j[�[s�d��#݉�V�5�ݯm��D��b�	�I��BI���ҟ ��ג�o~������t�Շ����~���k�@��~\-���p��}B��9v��mHU�W|�][DZ�&i0���c���A$���Np�$N�XI�b@���8_b.o���w*AپD��2��O_��ν���	�p�J���C����*��ř�=������ݚ|�}�_'�j��	*b��9űY��6�W�<�pIp�I��DL��צ��0~Ag1�:D=��w
�"s.~�{{��.;���3/W��mд�1x����>��HUXJ&t��jˈ�]A���]���# _�n��j�ѬM�k.��؟5�EPI��uY��B�P������2 ����$ҞHqo��WFzN�E������K�.Q;��F�:���7-��MQ�7S��D��r�e��*s
U��%7���E�X��	�C(2����xL^�� 