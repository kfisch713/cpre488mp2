XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ίĔ B���M���G?���ӂ��m\�����[>9?�ۂ!�~�G��^%DB��t��g��2��ɍC�]lf-%ߒ��/W��XG�~�"��7��]UDM����{�)���Y��5D�ܡe��$���ɚP�=�����3fU4º[��mA�Ζ�.������m�[�W��%�ˣk2z�"H��؆e_��L��p��֟>���c.���������f���1�'� _�b'����y�ᡪ�Ҿ6�ɾ����W�+UM����i��Lc�Ϛ.z�^�6u�� W�F@%��O��a��a���b��ܳ�{�,%�H�	_Q��צ��?ӦB����0�P=�/�u���1� ¯��&��
%��(kTgVn�?�P��b��N����8�c]j�� �rB��ŇCvٴ�"Dw��.�1)���g��4X��6{���l�&)0��j������Zk���o2YW��e�)��-��4)yqvL9��`Hj�B�9����H*Z�W+�d��Q�����ی��Y�N~;�g�vbɖ����7�&.��gu1�ɷ庩}j�_I%�!�&� 8(����7s�J\�l�V�I:R�D���|}��[9��n���_�ή��)E�
��!��I�A䏟q�Y��OЌ*�FWN�N�F�5�m)m��@� �Y:��LqTߺ��:�D>�!��y�N/�'QG><F�>sm�e���#�ϻQ�t��f�M�n�Y����1�:�֚w�`rɖ����֒EH���XlxVHYEB    fa00    26e0b��eS3&��ݏ$sԈ��jp�9oŗY�ikdLEʶ�XVА��W�1v��	��t�x0[#��/�t-�b��H�$3[�<�hT���(�A�4RW��~!��P�%�%�`*�{dR������-�`������#����Q̵2�anTyak�j���E��R�ˋ�����~]l���զ�K��*C�D��[Ri��£l�:E�YP�h�e�8����i�8�78dӝκ��w���!�A�A҆��pZ�a9���#�f*b�0�o��X;����	������lFcn�_�<� !S�F6 9�E��S�t���^�G�1�%=�� t��yG��-
�e�u���
��hsK�c����%>���f�R�T/�SK��`���'�y6�:�g�����(�ԒH�q�:_ȜS���^Z1�BG�������� �X�d��s5�[���P'�UO��=b����o����fF���{���7|��l��%����x�qN�)���=W�#9�5-����D��e#ôN��²mcKXt� ��N��x�lS����K�������A\��=��e}�x F���&U����G������ю�G����@���w���Q0�$�p�W)N�" �+���[_sC�8��U|A��/���ũ�>���`�"�,&�(�\�����2V������I����{)ok�|}o�>��8X��]nY%�͉r�4 >|Qeʛ(U)ƨ����!q�){g��GF�jY}�ÿ�!�U��PWQ��wB���|QrLo�q
3�_܌���R��Q��aC̊��}�=o �ޚ��}V��u�!g���Yث�i�rP��P�+*GÚ�V�N~}o�p��Y�<�R冿M]l`n��#v�6�Cqd�����ٜ�s�ad���5R5Y�c��������A�����S�	�t�?�x�Glt2��4�JH��!�\���\*k17�N�a�^��Կ� x<`��FnVq���>��N���6�`s����0����"���!���۹|k��0r�f�[=�d�g�3!�?�428���X�9���w"������e6����hu_|��m���;1^�1w���&����&Y�$��k�>8��ox;�:!ф�����Ͱ���{����|4���z%R��&1�4��߀��-%� ��g@?(f��Z	���6�������; ���{�� �XKb�v��=��+�(�	1���$\r�:Okb�Wՠ�����k�'Χ����?���Q�.I��>ᓖ�{c�Q=�C�@�-:�X=ǣ;vܾJ�.'�Y`��\�$�p��Dp��:� �G��ο�e)u	b��.���'	�c6-٧���+0N:	]�#Y��C��s�T�:m1����Lw/ �}OUM��GD�I�#�H ��	=�5IRˏ:�+�m83��6c���[6KuSys�ʈD?
���~6�sj��G���@�z'5/�Y%��R8��ga�E�-DY�T����}�(δ��q���*����(�l��JD�r���R���V��.D����@��>=�/.�����Q�٥����c�?��WE����Q�z�����-��(�?Y�1D�l�SM�Br�=H�Y����Fn�q{Ik�~�8	K�Km�ZNԚ�1�1��3�>���X6M��U*n�ҥ������*�l7l>ƍu �����F��s5�(����I;�ư%ϲ�2�r�
~�y. ���ܼ�T,`�I%ul�p��a��PVA���nϻ1�g�+��\'(�tm���UXW+�$��0����ҳĐ����Kd�>��a�k�6N�V@��bn�����`B�v��>kR"�Q�,R(����OA�PD0�gI���T�A��\
�o�ԕtpXٗ��@�Y�ӯu�x&.*�n������yR�0(
�x]_i(��wl�qO���5$2�Z�r?���办��n��7	�+/�Q� R�&�eO�;�'O�m��I8���d��)J����K�;B�O����2(H:L��!��*=�UwH1�ۛN�GP*,0����c\J���>�����Q8ڮ5�Ҧ�@:G50�s������e�*�$�F�N�F�rM���ǧ���S,T2�iz1~lZ��R���~�=�u��a�/��WJW���g�fو��,"SN0��� �?w��D��w��k���Y���6����|?c9�[�����Zd#a�MB9Ԡ��)SF��9G���X����뒾�ؾ~JL�9�aM�_h�U�I�*͂9Gԧ�6��p��������˻m]̦23�t+����C/�����ٻ�(+h1,8ҳN�Uh�%�
@�V5�
�{��/�4�'�{I���9��}r$���!�8pA���5Ƃ����g��sYM��M,g��~i� q����L�z8�!�(w�{�i�Y�'�,���M2%�/w�\��GO��/8~���$ƥ�"�\(����_B�T�ߢ$:���4��=�JG=q���:��GC��ir%���|�e���H���t0�$�ˈk=n�*N΄I�t�(��1�(]�+[Ad�$H�� ˾\&+�9�
1�r�|�����p���E�>z���!�l�a�k��D�ْ=oP�ω����ӹ}�U��$�{���+�����r�~m[�R�}~W٪���>!xu����9(�pK���fW U�)�z#~a��������Ce�g2��9n0 ����	����24��JG�81@aƎe���c<O"B�{���6���,�D��(y�Ny�;i�8����PDpP���9�U�T,��_U�^�cPXS,X�z�<����'�S����`�?���*1�ܷ�9���yex{��ۃ|O��GZ�߅���əy0�k{�� I7���8]��,��G�P�����!#��a�`��>:�NW��w�'e �����d?��?n2��(�1Q�$���x���fj}�O{��C��u����j4���%�SջN/�S����5x��a�.�L���M�8�:����PzȒK+��DXf��Q�O}m԰f����Ԯ4i,�mBg0&b�Z���m}?)MHJ�\�
�}��,�q��`T������lc��T2}�4h4Ψ���1�$:�<c0. ���@�Nb��g
(ŗ.U>��h����sA�R����M."F>�~�ڃn�;�:�]��&;p\�� ��@��zyăP��	��:�Z{�O0>��y�7W|���jd�>��K8��ʟ ���x}^�a��3s+>���1�.��Q�5�R��DCh��K�#օ/�x����A�\��A�����%�+�k26Ke( ���l{(C�<�� F���I1C�����~6'���/P�\�J�W6��O�Qgd��4KI����j�I/*2%R1h@_�t����_�O-}��~W2yX�=̠�ߨW�ᰠ�6 O�X���qH��u�0{��C����M�B+�র��O��3@�c'��0VZ4��_�4��"�D�B�ϓ����ѭ�Q�B��������N���d�Αc�L��.9���������*��l0�}?��ij���,W��(��I�%[\�>���*���=���8.�d�f���d��\�wp�ч���̪CX�;C�j'�c��7V�	�J`|�w��(��JQ0NY���U.��T��fS��
�$j�@Эui���O�3��5G�8�8o+{[�B#;�|6ߩx���}*���6d��G	�}���}����
�v�r\d#�`�x�,O�v�v���Xrw���ӗ�[sJE+�m��p#��� ���.b87+�}�٘�x�Wil�ESaJբ��6��0*S*�=��H����V�&��@��|(�x�L�3�\��<xf[�D���(M��~�f��Ѡ����g<ӥ��D�̪.)�d.�qL��,��c�o�9\�$��4G  ����\�'��"�]���H���4�Igֲ�%(i��kx�Xِ+��һHo�ڔ�u��p�����}��#t�\���� �KKH\[G'`ˬ�o�,�z '�n�C|6�O\&p|h3����S_�}���X�pb��s
����L}��A��z�I���[���)�$!+e��'e�\������,n��5c߶���^:'��k��["��,x�ֿϸ�>Br:��.n��c��u:4P�k��~�����=p%ͳGr��;~g@k6�Q��wV� 2�=�ۏ����W�!fr�g���ĵ�דB���ݤ�!��)tԙ [L�e}�?��ˢ}�O�6��9��xQUe�m-�a����|�?ED���Oea!9�?�R��RƱ�e����C�˶MK�G�Q��Ȱ���vNsyx��0��n�(�ɒvqY=-��Zb��K,z��]���AMƅE�i�f?���]�޹Y�A�+�x�������)����O�>�����:�«��h
!�øc&/V,8���g���n��<l�d��k�VA�)�C�� <p�qvV,9%�s�)(��L��ꠙ���r��<�>s]Uލ�����-�]���e�*s_�0��(�����IE�jC��[���F�i��1�t���X���S�,��l[VM����d%�)���Py�g(��۷ϕ��P�e�ł&�z����-��^T�%Ӝ�ty�U��ɨ����Zn��?  1<6�b�@��V��H�Z�5�|eV�>��b7{���d�l}�k<^�@+�����*�����"��nYm��[���v�+�0��� q�/�� �w=N�DZH��A^,͵������3�Ʒ
vW�8Z����;�JL�;ؚh��i���r7̻���ot�I~�e$�;�������_dO�/F�.�h�Y|�@!'݉�k.y�����Uո]U�w��� ��v�T5�l��T����((s����X�&0޾|�T�HL#`�\�ves�A3];*QM�� 2}�R��b5�i,B-�GS%Iy63�^Zb���"��y,ջs��$��3ʉbv�����oO�>� ��N��bD >?�x���=l�����2��.�5t,�>��q�Ӗ
H����pnQ�e	T�@�����Ɩ�x��l8�q�kV�Ì��� -$U#L���_8Nc���Z�N�[���{Rtܱ�S�*~hT��NNF��:��Ֆ�M@'Sη-Pq��5'�g�L+-�hjyLz@��ט��w���3��q��#�_�'�<F�Cǿ�b����#.[���3ιFH.J��᫷h�[�*��#��Ѕ��P%$��N�����j����+U���F���f�J���C�'L�VE���V"�2��3�b��� ��p-�L�)��o�ʼPxUdd���yX\/K>��3��@g�׼��T��'��-��h��OZ�&*Q�
ҵ��ry瑶Ϊ	@d$j��ȼP?ej���{�Cэ�+<9ְ.�e�˞ߞ�dqٔ��b�2���`�6��d��� 7��-�`m����ϣ�s���J��>#'� <��V!MI�]�|̡C���9T�k�g�	�Nn���A����u:�sAQ�_�
IN�a��cm�%�5��������"ݜyS�%�*V�2�k�pL, �(�f��M���1�oeX+|�]3�̖7v#"l�ܿ�<0�)\� t�D
2%@+0�j�ʘg�2��
��n���V#�����y$~Ԯo.1>�mN���SH��p�LT���5�6�����s.p�|�cm��xn
��"�+A��`ׇ<?U�,پe(����I����1��G8�)_�N��}j��~��a�������7�
{�ڭ�u�� (��3���b~��F�\��Q�3;�Sh�{M�tj�����ݖ
\��6W�T��-��z��=�:� ��^ܽ��}�Kt�m}�� ƻ�f_զKM���SY�U�+nLӎ���s�{_�)Q��|AG=�z�m�ڠ��=+e��3�Q���A��	Ӓ֍���^#slge[��!~Z�B�v�_��2jX�S�����*w��i��O��D�ࡘ�鞳a�$�����{�~ku�j_A��2Q+m>o�H/w�Y�l��D/�6���U��v��+�1,1j}�Y��=JN��tU��o�)H��9�kZ�������.��#���2��Mt�+R�ST�L�]er�2!A�5���< �����o��R[�<��'�Q#��z�:E�&B&?�5��'��_�fJ���Y�0���޴|UN���7��\��Pj�f�a�p�eXN��>�kk�^e{�Kvu��1�]&[+���tY�H.}4pt�����M�����G�O��ߜ��0��9��5Z�=�E���B��+ƚ�m�Z��%r���1��w��/�a�py�~�@�[���3��+:w	���>�6�LF�Ty1�ې�D��*�e1 p�u',��$�fA��	�;���	5K����+l�̂*��rB橬ٖR7~y��O�-6�PrV����됧�`����A�����MU���Fu�x�r�ֹ@��%�� A�T��&[��\�<��k��M�}_�eR'� P(j�j�		�l�Ȑ�9�8��7��L�V2�hB*�"�(qm�)�}�^K���<�R�*�jWd�6�2$Z��f�2�K�d��~��J����)�hS͊�T�1!}�Ҋ�*JB;�'�/�I��^�Y_��2*����@�~7�������ɱS�HD�r��ԣ}9�Hj��!V7/���i�׾�AQRXhK��hw�����bbw�aOZ�r��_����!w[�x|%�'�~��|�n��3R�Z,
�h�_�O�X�`��o����tZt����ގ>X��ޤ���m�BP��*������FK�#իL���g^�(��.桪�þ�z��^|�	@�hcq������� �_�QۍaChA ]��Q$�*�����U�{��a~6��Y�?o����^�+5�"a�f䝳��fԘ�_
J}Z�0����c��0�����W߇Y�$�|PJVK�������p��Qc�{v����ꒌ�������:�޳2>��qX?��d��i���$��p�
?�yp���i��fW�odg��2��T�x���
�a'��8@KA�(fK"��MT�\:!���읜��&�r����Aa���ms�r¦"����	`D/�c���,��������ͺ�������Dq�����y	�㘻8i�)�l��p��II��W8�zB�V��&�12���?��l��� 5���+!�SĮ�N��(�oxg��ʿḊ�Ө�v@0IZ��+D�P�z��ה���s�]�ut��8j�}^�$-�]����L�MΈ�(�(�Uh���L�"E��F�t嶆����!�U��X��G��T:�$z��zʕ�TGĢ�c�^A_n![-���ɫ��+bM��T�j!�F���eL����k����\��3?��/���?I��H�&Xk�H�p���%��udrG2f��S��=J2.�q������� ��7�j��v��ƒg.�m;����m��v�@�jb�I�mL�K&�Xk���P����-D����._ɨ���A�A���z�G��۠�ς>����.���zj����f��]�$�a��W�G�~s�rB:�"t�ě�Z����^��%g鸲2y��H:iu/�����3/�[�J��������,s����,��yPKd��o��bZ�0�R��,V�Չ�=l	~pK��ER0�w;�5L_�Øp���ex�IE^1���4pnXY�`��S��`��t7����W�0/�/����!^���Ë�}�3�H�c�3&B����4D��.��\\[X�C��S߽b�fD;Bzj�ó�J� �7�=F3������	�@q��Y}j�WTeCT}�k�`�8�܌�L+�o�Z�������v+I��hY�b�ė�jJ��0ِ��s�nr~�WX�|N��X�:ރ��Ta"�)�p�9�)W��!��[���N��Pך ��wlO^�ԚL)1;r��ʸ�2m�2:��!�ce���;��+!o얀�_��������gn��tQZFk����h��n�Q�F�2�n'���V �TKe�8ZVd BHU��`h4u����Ċ��JX�� W��?�ϛ�`f�Ӗ�,�n�g����ԫ����wڢ+�`N� n�T:�x�} \ib+�~�lO��Va�C���1��_.�I!ҫ��:#j!�_���:�}ߕ�1��hu1��\p&��Ag�??�:(�7z��<G@�rG��1J׌a��Fl�7�R�>�˙Y���`Q7�� ��������Uk�h	P��PKϐD���(�?��'��h����~�
���l3͔e1���i��cܭ� �SK�[\��=Z�P�iJ{���(]��S�~C`�p����5L|�?��������]��OL��5B؄�m�H�����O�>�9:
t�Ou0�?B�2�]@���_�F����l��0�c`l�JJ��B�)������ ����r�5�$u�0�?����h���-s�݁+\
1ok��.��6I\"(2�RD�X�Xށc�r�T�ߧ���ªՂ$7�������� QS��!JJ�+nl�z�1�r��*]/��@o^�%5:yXc"�ɼ=��L�=�:��\#iz�Q��Z��C/쿓J�R{RHn�����ڝs�u�Rd�k�g�Vv	����C���+U������{��E�u�ų �X��)��CI�FWF�V�DE0>��}�Q�燖�ZW�0� �s`����0�9R�aL����L�������Ru��_�y�#6�jT	�V"@9��q�6�{��i�R�^�����*������/��Y<����x{��B��6y���uV/g�<GN���8���?�3*:�%��x���/��2{%�5��e�P�,
)���s@��X���.�������,�7���������u��a��F@��n����fwe�0�4���l���0/�6��u�8Nx�60�jJ�@gt�5y�-�[�TE�7���X��%��>���%��?�Q+�RLK$� )CO|~��*��h���o�+��heL���R/�yNz��W;o	W����p!�&'�)�^�.�)A
��/�1�l+�M4�z�S�C�o�Ć9�7�`x
��+����xC5�֔'��kh�����f����RV���^��nF����F����P��pk-�\����bm
�ɺ+��fI�8�N{_�&ő�9u��D�OY=X��f%�4g~�	�����:"_�)�w�#D��y�D�"3"��l�?�pN]�������i]�
8���rcљ`�	s2�g��]NqpX���:xn��j��=Rh})����YL������<�}.�k�;C0E'��m�p�l� 
D&K����\:���� "?=��j�n�59����B��� ���O���@Qb�o���M�.[|��F��e���������`Š��_��8�RD��t�9"�*��� �ƚ�G<���+m�U� V��׋��	"�GWR �9I<��|7��YɈ_�)��G�862OJ{���|C�vu�Rc� �%( ��ӷmi���	c4FpU�C��oO�����9@$�Ū�%�c��z�@���* ���$y�Zp���}X��rX�'0�nfr/��#L(���8�����p�XlxVHYEB    7d55    1450���s��V�g�t5��On���"�+b@&����dzg����>��xP<$�e��-xI����=/U��	�XJX��g_��-�]@-������呢 �-���__�~.-�<�L�M���@j�Cs��	6�hH�.RR4h�W��T �|�-���lï�=���4�T5L���N���(�������9��+����)B�]|M�^r�D��Ƭ��=~-P�vT���Nw����%��mLG>J�J�J�p�4�.�_O�_9Y��u+W�_���1��8r�%��!~A�(��,��r0���σSpM�����_�Vr�3��w ����?:�	�����}�n������VE��w(	������K��ϧ|B�d�����K"0���v�4��M�i=����N�=�Q��Ǹ��4ZUL˻�sqgROta�FW��Pt߽ݼV���ΩO\�"I�jM�gtqf�#zT�x¡���2�XI7(優E���ZM�Ά^u,L|;���]n�Jolw7FX�jMbv��T�y�%�A���ߢ U�: >k5�T�8���Bm��}U�[����O��V�X����4�������)wu'�o\��4���wf���J2��F�@�]����5��Ԣ�o.>�e�Oc9U�GCN�4�r{��
l;�Z,InL�.��-Rt��%&��%GQ����4ߞ�,�`�_��|t��ɛ�P��m�&d���;��
�Ҳ�p}�es�[��ȒJ��;�w�q�b�e�e�g����@�pS�{,���󔉪_M�,H�e�f'��R�55�#(�jD�_��\�����[c[�)Du)��Kc_U�O�$
K�Ms��wT`ȕ�ʪ����\{�-�6m5+��Z�Q
C���Mȑ�M"��[T{-��ҥ�`�S����YQ;��]{���L�S.�>aװ�
��>��Tx	�7Ӹ5�����#Q��e���3�Uȏ�܍}QB�V�K�DAy��с�-���[�0�pX$��m�c3�g�^��QL�ZH�Q�N���<UA��5�̲"/1ͩG/���bV̈́��h@]��!S@7
��^!���SJ$�~�R�#i��el�*��޷�w�G���4�ח�rֶ��}��z� 6��ں��M{��g�6�|�xDsX���z~[x9vq��V�\u��|��N�1T����;2��� ��7ь�M#+�$X�LQ��9��Zf�}�3�x����a�T���u���{\yڀXS���=xW�e�Z�+ļS�p�I�	l�w~�Z�93.[^�䤁�#��qr�b�V/��O뤷 �dY�{�z�N5��*1����=:h�{�.BR��h�����R��ͿJ@�m��M�gH�\ιP�vGЇy7}�g*�}�;e�.���ۖw��~�s������)u	��=���9�S���ÿX��)�bfl���m c��i_���G�$����'Z|��Đ��+�Q�*:�L�8���ţ� �;|9����F��ί&bx9����=a����F�H�q�JL�"����}�38�����R��01��O|������+�MAh��� ��e���8_�#�3�&�{5�}_	3{T�����`N�43�'����ݮ�$����~d֫L���mp�LC���bbHM[���w�ה��ق]GHB�_67����0��xRu�[�c�w��*�����NƗ�%�+A��yTr�����C4�����(�����̇� ��"K���e�'�i��~/��,'��E?!��>:��Y�6�|M��@h��n��c����X2��_���f�ł��Y��S�>�;��;#�U��|�AzV�a/�$l�2���vA�D5�'&�-�I
���ʵ+����n*�,�z|q�Q'�ӒB�#<S�u��.����[uF�2�
��j �)�����~S��bɯb�e�V�4v���������Rf����% �T���o�G'Z����7x7�2ma���DͲg�����������nRDM�8 ��$�6o����o�Z���%{�eY���cs�O�k�.����6�F�,��fi������wD��=/U����2�t��&�ߚW��<^F��e3�u]�c�a�q�a\3En�t��k��g���mq��XM���$�îcl�'�8.d�`���� L�E�S9�cD�Uո5za�1ѓ9��l��`���m��������G
 �A�3��V���z�����/w�Ŋ�N�/*���&hA�;��k,w{�m2�]��F�ݛ�R����F��$�V]Bcu_�
�;�т4 %u���~�g'.&��Oڢ>>�fG�_��w�j��8�������u�H5皺�y�(�j)o�?z핑�&����� ��f࢐[]��=rBP:����s)W��N�7��xv��]�x�B�ف��N+��n2T@8��'�XE�L�T��Dbyn;*`M���&A����р��Fع��N������FI>LQ�M���tn����+���Gy ���x_��{�6��C����?�Y�6�+6���{�z(A�gL�����#��c������1�>�|#���K��W�n�i��9�g=ŉ�i��V��r��s�����t�:UM�j+ec����{�/B8��>�\S)ʜ�Kj��a�0���gΥ���&�[ ��X�ضx��)}�2)I�H��6�����b�i�%섗�~�Y`�� �{�]��ω�F�R	�){f�����i�}��
0��hF��ѣCmϹ�^�e�vgb���f����L��>~��xY��m�m��z9�3����b���;��)'�����cA�������' e��rE�A��/�I��������c�D�Vc��7��زCL�z��vF�����K�ꁀ����d
@�Z2�\'���$`m`��-��O�?��HSvV̸���FMW�(!gn �q�0�V��%�#q{��>d��*��9Rx�~�u>:��TGƙ$��1n�$*�
F��`���(�䀦�>��*8�
�D`����)���I�����'��g�����-��1�.�<��S�np�L�F�2�|�zB��.|Dl�V�R��8��nD��̙݊��I��7��B��]�$�vW���]���aB���!�M��d�}gf�N��ͷM�F��������"혲. ǀ��Ts1�h�8N,6�BT8$����4om�>h��i�L�N�n�����˰�s.���7O�#�~B�:���&nVH�EO6��S�߈'�Hhk��A4��r���!(ݘ��Z�rFv�uy��H�*�5��7V��wR��ϑA�I�r���;���7�HP�<�"�������B�b��������䭓L�c񉈽c4X�^���mf�վ*g�����A��?�٩�"\��v�i�em��X�̬4E5dP<m�Z�r�T���.b��kq��Nx����u�2��o�WR�.~S�<}�<�!94l�Fk��d�屠�Z6=^~���=�I𢮠|N,���!B�_zS��
�sF����t�Z�@C#ʽ����m�/D���>�tA�〮�W'��&��@���eA�|H
��*��m�OEv��4g5F�w�Z3�U�ǚ��E�����G|�C�Ne��^��S���!���x��.��ǲe��w2�?���gK��O	�wk�K�)~ZT���y�6M����*�Y�|�4k�oQafK[r��%�J�*�e�����l �{��:�ޡ���Eʆ�ߠJ�<��V��GI�F/�a��@7��-w��9	��B������iDڌ�`�B�>�u�-h��
>lU�oASe6�.�ª!�3��b��_��:�n��u)ߎ�W����9�E��u��`���y	�q"�ؾ�zrK���X���"�O���E���L��i��pM�97u xY��$"������s���jL��Ց�xِ,x]��:K8q-
W����G�z̴%�v�.�Q�K�<��J�
����'�ՠ?��?.��C:G�N�������')��8�r�N��������M���A�&qq̵,g��n�?�*h�p��|ɧm$b��}���-�ژ���X�ɕ��`�.���z�t˷&��v����"فq��H!�g)�G���O�y�j�]MO�Hc��H�ͮ���?⣱C	��<1��dG}���G�e�mX���v��;Q��;D��JR1R yᎱ�$:��+,{�{� #Ă:�?��*,�B��|��MA �h;?��'�x�ݔ�l��E�> Ư~�#���*�P�[dv}�)���9<�oi�RZ+�#@�]�\���> F��<҂�b�4�<�,��/�^�t�)�է��y�������� �&ۙT����?���k���N ��Cdʈ�.�����\�����-�0��>��{L ?Z��Pd�Jq�^R�k�bp�g{`�}�hO؋�� ��Ib�2*Ԁ�����q-��i �H��rW�����:���]XP=b�O�G�H�+�g5SyYt�h�o�>4��9�3������z�Bk*��T�L�Ƈeȋ�=br�(��5����̥����op4� 
��i�����[:��SB�{�g4�>u��O��v�B�����C��*q�$�Ph��=XI	��7J
�#�!�R�DR�Sp<,��kvA��;�<5�쇍U�τ�uR]�<���¬=�X��U%�#�%A��Kk�h�vO#n�^xM7�Ba��`���Н�������	sjk[���Je:���2�p+�#Y���S8 !��L�HFE�Z3K�* U��+�`���8-z=&~��
v�H�y����h�v�'�^a�ak��ˈ%c�m��CQ6����n�ɟ9�a�К��n$���y?�4���e��	k2V��I9�>�:4�wyi��KY�+ih��������:��g�n��@��R�ǥT�	 h�Ҵ�Ő�7��K�N~��9�ۧ��\跒3q�*�`]uj��R���]7n�_D��G��L�W�w�+I��