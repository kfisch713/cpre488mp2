XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|#�$A�ԑy��v4Bו~Q�o8�^~C���|~B�lC�����S�*l�m�B�<�^��"�_���5�/��#�l�7�E��T2\-o�����XJcFnP��h�J:>��?�����2ܜ":o����
hoP=4G�!� {ښ�����l���s�<k���X�ȹ
2��5�Q �Z���?�oF3p,�00gU�49��c�k����Zď�-�+(�8��迴
�N�K��#�]���G3���ϩZD_�1ؒ��B%̔�M7�{��ʧ�^�R�}G:=`G�(0�@Z%����G���U�u>v��h�f՟ h�1�<�g)a�Tz�^o`0�!�D)g�,9��?mckN�yS]���X�/�X?(�Ŧ��T��^�\踃��m�ê��R������Ք�r���-�6��ct/_�a2<I��Ђ}���z��%p�P�B"��Kwrwm�]k�~bW�c�t��.K�JG��*��f�
 -��$c��j���^8�E�T�ɦ���5H���4I��ghMEI*L1s_��)�8�<�̔W]0dҖ���QĿY����֚BE7 �.����S&�-����P%(��k���2���H����a�JE��QDe�Ѩ8~��'?�Q=S��b�d�co�a!Ĭ�SÓ�\�*o�!��O�6��!��F�%�e�$��m��g��]YYС�%��������a���Π�(�>�]:��2����.��T��&�#�Ù��ߔ^��D�&1F����f8p�Q�ݓ�XlxVHYEB    290e     af0BE^��|��̇p|�(��7�}V�Ҹ'��ZS�7�]�����3|�c���q���S�lĳ��w������f8��%�����s��~c�]ڣ�%���v.�������J����)Y�X��OR�c�C ��䡾�^-P���m��&�oݻ�L�iԇ���QU���wI��]�kJ�1#P�T�U�v��W4���0�����p�.��������E�-�������b
)'w0�~Z�����������/9���6�G}��jF�� j����w�Fګ����膛p���/����~e�6�j��S1s�8)o�
��H�Ѩ��X�4�*bx�����<P޴����~��7Y{�æ�>]����r�r�n�G�'��
v��P~x�,�M#<x!�T���AO�ۖ�[��蒬�8d�I�OX���G}Mb͜����d�3#E)�j�S�g�}�!�����=�T��*�g͔n�zV)�PU:�TGob�aJ�sī1i9�O�_* �������ڌGh���q������Vt%����+˷B!t�} ��K!%�2[;�CҦ.�����;�;�D'�lg���)�7����}pٱ�z��A�د��GB�]�\���K�� ,�U��9OW(c,U��{D��N���k��L}0�%NV��e'e*1tf׏����ol������M*���g��N����n��$��x�1��ÕpI��3N׉�m����,?aL��?��
L ����l��,��}���[�d�,g3�۫ﵮ��q��q��K�熈���~σe�7���.�N�<�������\T,�|���č�g9��M�"W=��g	����";�ΡT��f��Θ��B�cQ+g,�\�N��ۻ#l�nv&�X�}�zi�0A&�/_;�t^�Ю0�9���_��S���{�yT8�Wbb�I�:�ZS0���h��r������3�f��[�N���XV���W�v������P�>n�
M�Z^����mw�'��h�ܤ�͜9�e��5!����3Sat/�Φ�asg�#��A1���A ��i��R�B������/)����E4����ː�����0t��?5Z�@����K��V5�j]̙MeBS�=��.�!�}{�kU1�H��s��:��t�9$��(��)���%:W��l3S�y�"h�*��Ew�C�BC�H'z�#�$�[��cR
xq�0��n�Y��1�z�ѓ����L4��lx�RL�$z�i�'i��qg�@iS��*uBh)�*��9�<QE'J��4��*Қ�f��d�Y������([����(�D��H�p����D�-q�U2$`I���,�(���o%Bcan���013zae��E���ܩ�|Ka�ش��8�e����f@U��yO�y��ה��5q@��KQ��tE���ѻ�̜z������7j��q�nH3�cCN6Z`[D`A�w�?p-�`���nj���q2 �:��aR&���
�s�t�Y����ӈ��_��R3����#M�Xo���~Z����R}8�8_�%�}[����57�.��o�gr�O�i�&G�<�C�w��8Fe>�A�9A���2)�\fTH�]�F����� ��Q����By�%SB��$��@��D`� fs�&K�8ⵘ���L��Hv*`}7&v�G>;U���Vu��M�Z�W�0r_Fԁ'M ��e�#~�g�a� #�=M�ŧ���P+ �*��)�j7.�Њ���-.�j�u}VBm�o�g�����{RݔG���)I|�&�B� �+I���!�"(*�O�(?_Ё��H���[�?���_j����s2�JJ��N��2֙���9��%�Z�%b+����:�&��Ė�����е���8�P#����m|L�L�M��֮�2Ø&�<~�؍Q��=��;H��qB�ܦޝE�C��9�HeG��\_��S>گ�'�ˊ��N~b؏Y�X�c�*����L�����-
���Z�e\���h���})C�lt%�vE��QxŮ�joQ^N�o�=�/]��%fY���ﯷ} �m�#ُ6�D'�����z�wb0~���-���Ơ��	 ۥd�r1)�Ǜx�ӵ��Z�W,�ِc��d��4��R���w}�̗Ԟ40fܲvp���N�����:���"H��u����t�z�{ca"L��&�%$���:M�s۩�P��N).uݦ1�?�i�ԜmHCeM]vū�]���u�W�:-!c�a�ֻl��Ŭ���~�z&�96+(W�X�]�{���ϯ�p��c� �y�V�����9�U\x�YvR��P�q��tyL��1�=#�AT��Ɨ�k�t�S�v۬��l��j/|���,_�Ȣ���v.��k�ɑR4�X�C~�v���P��"���g�ۢ)c�t0�w�%2��G��1$D�@�0#[.��Ya�N��TSQ�=z9���z�u���������L8�Kz��ZU�)�oy%��؃�[�&��괬�nl���.==T�����<I�8����ސ0�E�w���2�1�DY�F:�FA�ѥ��괧�}�����p_�}�Xl�7�r�Cmv�ρh�A����8u�O�o^���у��)��!�9����r;���γ�Ew�A�]�5����uHr栚�Yoyi*^���%�~�RϽT���Z������Vb�3�(m��g��rl����K��)���U������Hg�qm�u�hN5���g8