XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m�#U�e���Ґ���T���lb���-c�@�tȢ�@jMe�֦�;�7l����8�����L��чk\�����=��=Ǧ�MZ�Ԩp�'�����n�V�d�#��P��S���O���D����/B�8N��� ����rvY�B������vp7������F�ԗ~F�������{x(��2xzY�~�9ځ�L�Zƻ$]
_���su��P�Dt���аv���'���"�^u1������P�՟duQ]�~�uc�*�"�M�*�]��5F�9��VP���}բ�D0��b �������|��l�nv���?yl����Z��|`"ť)���֞`�iwHDӻI��]�{���},��hNT��Q6t�ՔO[pZg�m��:s�q~�g%�f���O�˛��c��7�$�|�/���m������Iu�J�_�zb����L�S�^�.)�я��,Q���"���1!���� ��>��՛n q��̱T� :��h��Q<Z�"#��v2z�6BӪ���f�&��qC��CU��i� �,�R~!]V́�>ᾛ�5�E�fu���g��xQ���f�����F�y�'C֯����M����ו5��5��t���F�$���[�펑�A7��eeEl���H�����H8r&o%z����}nE;)���	L?�Y	�j�����GZ�n{5�@��T�\��;��$�8��#c��6�������W�m�3-;i;a$��3XlxVHYEB    5866    1100��
�Z��_����T��ѥǋ_�|䝈)o�0vΔ��}S9����2��b�2��J��D	'���R�m���#/�JQ��7�vn���O,i3L��&��I"��dZ�g�sk���<��L'Q?*�	�R�Ha;{�@v��ej�t	=31�-�O�����l�����r֊oW�".�X�ͯe��{��G��q�=ϠcV��HM���+X�D�$H�x�]\���_qe����T���?�P!�GڢY�j� pN��0U�[�>�i����-\�kBc�r5��כ��<��x����U��j{��a�����T�6+&/���g-Ў��L�j�]���)�pѢ6�0�XZ��lۢ�7��`f�>͵��?(�@·L����z�,s���P�� ~�Z�g��'[^̢ S�*9�"HeU�+��)+��ٞ�� �F���6J���k���8�R_�{l���M��M�l��(�p7G36/k���(}�;��vpZ��Vkc�MΞ�[%�;���/h 4�UG��;R5�P(�G^^���)��3��e����Kc��q�Sa�%���Lyy�^]�܍�-��x��?��mf�T�{�IFshE�nP��;햼/�@��ܷ)����#�)�� ���~u;{�I�b3��uE]0k�A`���`�8Bߋ�8Oρa���Ԅy�5�Ǟ[&~��k�Ԟ�z�w�#^��G�x0�&Q��V�Lji;ei�Z�r��< [&��6P��N�k���-�y����:��ϲ~��:���<�26��yw4a�2�I�~�n���W�o0�v"qSG��>'X!S�BY}��U�ݤ
4�8����
T�a%����P~灺��q�K˰!�sɸ!��V,�������GĳF�N0�P��f�� p�]�l��A6���X'��T�}h����\B�*�;
B���a�]��~�H����T'=b������N����Q�� ́T��L�?g�5�3��<�y׊μ������s�����f�
��!��F�@1�ܬ)�	���X�@I�ǚp*��`R�����)p/&��K�ZF�@u�]��[�F!���@���ϊǑ�7`(�=L^s���uR���(��\bB�p���)f0�&��o�	?�W�ܖ�f� �P=2
�!ͻwk���Wv��e���2�"N�?`�ȦIT%"0��	��_+�Qr�=��Չ�HU�k�Xޱ�ۈ���Ÿ�݆��2g:�� ��_HL�#��z��,���=k}�T��� �ʐ�,HZk13�c��9���m���tv�e8���þO�o�(ǒ���^=vm�ivV�`)]�!'1�ފu�z�lrk�� ���I��y�M�b���N�b}�"	���e?O%E���E��	��<�S�"�l/����B����U�b���)O��A:�7���s-�4���R(�t���8��rTU���a�Ԯ!�v `��q����R⿥�wc��ZP92��.r�.��� xI��������Ώ�$����Yi��,=�<R�Et!�X�oť4���-��zi��h���8�[�D.��2�UZ;��t!Mt��a�6�q]��e���^��D��x��v����.GƜ��|1��h�|}ŕ����X�n�XU�G�7Q�u���8Z�Fn�\����Y F��b�����]���B���C��g�_�OP5� ��q��=��z%^��	U�ͽ�s;����0�4�PUZ���2���z�a,�QuV�O��a�C<�N�{w��B~��l�,(:��Ƹ6O�uɯ�<M��<��^!�6a�bj�������1��D��]_K��o�9�$��4\58��#�,�Xi��*�m]k��C��	p�o��(��"*6��\8�R؜���&w�q{�TC������"�:�l����LᬦF��&Z��y�ETQ'F�l��3��ҳ,����J�vϊy������L����2doNۗ�	˧b�����u<4�??��@i�_�-P˖��9>�Pa, P�ϤT��q�̲!���w#�f7��j�m����\��1 G�ti	�`_%�G�P�{/{�R�}��i���)�EjS�LH����$B�|��&3�rla�껛!!��b��#��_�4!�e�`�iF�	���Y� ��9��d]������X��g�����^��y����Guq��.��R�[I֡��+�q�b]�!NY��ba�S��(�}$7�ph�0��yr%!⢑�4��0����|Q8v�t��o�^GFX�A�e��j�u��+^�1��d��p��8��4yw���Wb�"V��҅�ԗ����A@�G)Ykݐ���D��2�.�ݻy�R����/��j�[;�wF�d�m�8q��_7���^� ]��a�~�d����0Q��V�(��-�Ifr}����y.�^E��K��fO!Z9مZ�5���D�[��I�1���&������H�U�IMHYC )����4P~o糮xqQ
�naK-2�nL��q}��|���Z�����D��V��2w�phZ�m�{�MG�\%c{�I������9��>Vj���[2P��K0/����V�	�Si�7
�7М:��QI�xTȉ1RH��ɗ%x�_��-rg�'��4^�F��CRo��|�&@wb~��	{��o����WΛK@ ʗ�H�x�ä��	B�H���%��T� ���������N�d��Z�Sqwi��)7z �K��@��Kܣ�A�ц�Z����0�'�(���]�:��XAdvXE��w���ب��q�m:4-�n\��X������q[���x|�S.�c~�t�u�a�����s��cqU��O�;�j�V���PA����0�8v5ެ�$�MG��O��rg�177�jc��%+|� 	�]<ϱ����r�{�/\Og �\7@������7�P��O��b��>9��>9�6�U��s��U������mh�����A����@�ˡI0�_^*f�y�h��!���:|��9���f$|�CaY����ډ�i�"2qvs據v��6�Ј��5�+�T1����y:~#P�t���d�JBQ<-�Z�cI���WF��'�t�tKGbK�e�?u�*�AS�@s:2RL�W���^�EPCm(Kx"l>l��V���b]ۑ��8��.�:����&���h��VF�|�Afe��L>�XI�kX��/��P��*,d:D���AQ�H ���X/I����Q|DI�;0�o���l�9P`/S47R�)�o�4��#���$s�*p���oXb �-��g��2+l�ŀ�.+%�5����M+�u�v�;�����[�:$%���(J��}�	=�p��������ʃy
B�~%2��D5��:o)R#�4}ޔ愞�:��&edo�V��\�=��ОY��k�
�\����3m�~N�a�<ޡh�_�;���X1|Y[�o}+o$��0'�n�v���P7��B�G���|iҶf�d�7(����r39�ܺĹ���C�U�Y�w��6�����;�d|�����)��Qݠ���u��s�c':��JGS�����$�hN����n�j�+@�G�$N�S�g<?[��3�amr�G��;�e����W����U{�<�Q���;�8��~�n��%#��	��V)� W��%4��|�rI���X\R����j�y-sk���3�s��.T𷌶���*���s�������0�,0	�14Cv*�����]�dm��\@�I9���'���
}T��D��F���Ҋrh�C�l`E#"��7{��*ݽ�X������#n��л�
� �9Is� �jP&N-�7�v*����_�F���f��6Y���������~�5�s��g�:�G�jy	����|�u�=an�J��y��ț���ƿ>H��"���{�'~�_r�\����T�*»z��m]�^���o��e-��
����1x�����F�B.�EL��n���b����	8�Q!hIb�3mQ��bԩ�Kh%:{E�h�_%)���6��/� q�4B~��(�t'��]�e��$/�U[v�"V�;�ݐj&S�@���8�xվˀ5�A���/м\�3���4꾚�\��B 3�����L�*v3 ��.�W��=���D���;�����]�(R9��=% 3��++l6vQ��mwr-���Eπ=��q(����O�@���>��bqD�T���I�c�&q��:�<ۚv���RI4}��Q7�r����<�d�T���'�_��U��@���