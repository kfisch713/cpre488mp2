XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ģ��,���rt5�V�%3-<0�>1�H�+w�s���'����b�K��?Z]���.�p0�W�i#u���߮*�Q6��:(�S���1��ȕ�����r��1��{���!����� �i�h��&����&H�(��b�O��d�y�����B�w�r	���wg�a�wU&�}�P�$��4����9�= V�4�;��sǰU��π�VE{w^8�n��ʱW����Z\�N}��{�S=�O���_�G���ֈz�F��Yp���p;5��u��L������ъ�5Ӏ�0[��(�{�I�l�~�)�\��h�=�K�B}Z����C����(�Y��:�I��_�]��^�
5�Aee�>ϐ�I@���`x�[����Q�L>6Y5��U�r`$��Iݔ�.x�{7|�3G��%���t�&2#������ѝ��7�7��/]��}f��n���N�pEʙ�GV�K�-^alx"��f%iZ�:a}u��D�+�K*#�|$���\�f{s�k���a��q_��Y�����g ���V�n�ϲ!���?��#���xsa.��B(�ut�e��� zͳN�$�]`�Q(�p�,�mE�e�=U�����2h3��<���?.���m�M�~`�1��
���y��U1k��A(Ȍ��TK&o&�����L��W��ع��8��̸Cg�s�*cf$�$��h��Є�W��Wvl��Ab	��4�$
g��XlxVHYEB    da59    2e30�~I�>�G�:S�ӢU����Ϗ���Q�IX���mrG<s�\?��c�H�����1���FG�;��b5U��;��X�Tю��Q��	�u��4'��2��n��rJ��sB���;9�
v�x&���`l4�.}nn�'����*�����yj��J
tM>ڶ2:ƒ�>�0��r�[���`��s=�z���������ko.���0�ѷ"��*%��E;���FC@���>��Cvy�BB���kw�Xg�Eوt�'�!��e6kg�>�E%�R��d�Bv�S��16ƥ�&�$72{�p��E�:��N��3������;K��%��P]
����߶+�"fJ�)�� C����-�8�ԐO��ݱ�W�����cFAIy
>w5H�ZRR����Z���ޯ��p�Cĥs'X�z'�M���ZA羉��|�>�Ř�P����0����(������U�����8[���d��f�~?N�Qk�7��4�u�ݜ�A0
�܀-�)LS��5�o��Z�;��q�$c�]��/B1/Bz���9����G�p���^����(�j��PL�j��9�	�+�[���i�{�Km͎[��&f�ӌ*�-_D�]_q�
ܼ�X�v�P�@�cb��չ�y�x�������S���؏�����/�(ݹ�o��ZU�{u_�c��ӗ��Eɶ�Gx�>-��̗�d(���?�~�F������:�����G��sa�a�uE�,�4)�۵ 8��_<�P(�����z�\��a�� 'ݯ�9��%F�|�*��DaC�����u-�#<��@��Ip�.">o<"k�:}�>�;�F�Q������ú�����f/���=��s������҉xN��5 I�?0�j�뫳��7����#mO�'�q�dW �����8wӵt�E\�Ďsi�+>��d�|�"�~9mV.��(8?�M%X�P�J�E�p�	�W5&�����+q�/tɗ<sp����*x�� r�;�sq'��ϐ�bI5�ce���T���E=�|7�ĺ��a�r�?�r����B�a�jղ�V�Y���ġ�o�)����C���Es>������3&zW8N��W-ȑ��@\�&�F�*�����?^���� ��U��!2sY^�ə��{�z!�p���H���26��㰩�� ���D�y >��N��X�"�yTߥI�z��b�H�� ��	��#)�\j��=��ѬXNg7(���.����P�� ��[@�W�}u�S5�T����=�h4n��q1l�un����>6�Ǫ&ɀ_�r�x(�`����xb�c����Nq���o�e�"hr-:7��@!w䮯��M��j��<�8otv�a}���/��v%s�]�C�!.�/�T�æٝp��1�u3V`Z�9�9]	���h�~��a����H3�E����
A�_E��(4]��f>fBTz���VT����b�cg��p�I*�J�\��#5�*_���ßD�3�x�#��)�h��������X�bv�u���=9��{4+�Q�;�W1�NE��y����i�3YfZ�s�M�+U9�$^��h�y��Qm=�틾4]e�����Y���nS[�x\T�ne����[OT���'�ܟg��`u��ٵj�،�f؝`F��s�@��]���M��r6�EHH��lNR<Ђ����'68_�`ֽ�N��{�'l����,�י������6IM���z���J�Q�b҇QV�ө����9���{/aa���2��mC�j�e��l�X�#��V����G��wQ����":�kC��j��q[	��]F�{���L��G�NA�O7�9<�W�vNg5�H���M�xvط�Y�
�}��w��>��.�S�3S���d{B^�@�y.��4�驪�t�����γ�)!3ߣ�q؁kTrW7i`)�����O(��bl�zS�g|WK���𓝁T�T���S�W4�5�aF!�*���b��#?N�_�2��8��
�n����]�4�	I�g��w8��v���ւ�o���E�Ȟ�:_z�j��umk��i��7��W��H�@B�z����l(�o��d$_U��[>3�^b�7e�;z�6�`��=�����:��.H��zmA�\���pDm{^\�]aD3��K�M�ES��"=0�N����~X\���:��˕��`5dÿ��I�Y[�����^p�i��j�8i�q�����lY�Lj�O	e����Eߑ�� 3)��&s:��&��j�Wa�qþnA��4> ��r�61����zt4=,'��ʼ&����M����$�V�O�|�oL�,�P�H�3�"�i��UVY�;�
�>Ln31 ��4�i��u2GR�eC��������'����'��v��;1 Cx���Ǧ��"��Ax���p��8m�C4�}x�1��~L]3�A|���6����C5�V1aְ2߲��?Xf�ox E�R|��a�sAsWnuX�w�3?�q?r�/[�4�w��C�[/��o�����v ��8�(��^,�8��7Ht�U[��_lM*Q���W�����"ceUp�ΨK�{�E���?˱B��?�I9�`��p��f%�TR=���c�k1��q�4ҧ-���=J8��t_G�R+Dſ�SD1��*!JN��\��7�њ�C����mM}n��@:��|�pհ�/�#�l�Nu�nyޗ���bU%���C����6� ��f1xҤ�*����-���-��|�,}���>*�!�jl��W�D�t��$��0B{��=��{*�f�I; .�,>��,�LU��Cס��"��rD�c��W��� 5����_��=jv���'�<��')$�X.�3��"����>�R�%�71�|ZNqq�Xx�&zi�/7*d!�V�r���kB�n�`�_%5?��v����.q�Hr|��J���4�&�0��R4r-c��>�^ܔB2��w�d���
^}�$������٣ًj�MG��-%lB��~����q���u�.^V�����BJ%�350q�yT!Qu��lL`�v�%���w�-_��J�3�]�x��xM�c�A"F��&}��>r��ӟ��8t�s�z�O�J��V�e����xOeIfB?���W!e&~!�"�y��k�\	�k2��UNm8q��OTT�#y\�|�>�MQ��>��%�]H�e$N��d�C�'��j��%���}ϳ�lfд�1���0N���a��k��MPTI�u��蓠O/UB�k�㵼�eE�&sQ�4��K �،�f�]A��vYuYny��a26ӣיʃ	�Ԣ�Y�U6h<�gL^ha��S�����`�@i��"Ѹ� iF������'�:���tܰ��^w��B�}̚�V�R�} �>� Ͻ�l�ɭd3���]x�~L�ap��
c�DK��5�ӂ��O�o�SԘ|I��]���j"?��W�Aa�ipEIR��8@x�:�p�RÄ�}\u��5���K�� bY�u����H�#o�>v	�{T7�N����Z�d�\60}tu�������0���)y��W��;aH�
�-�k�ݕ{�AR��-��(i�
�Zݽ���D�/ь*H��h�#��=���:�y�M֕$��O�(eo���C�9�y4�(�HQ4��҄Yb�S�z���X<��0��˿�lS{.>�^�w�آ�����a�_��N:��?�o��'T��ɬ>Ln-��=��8#�Ɂqi�/Ο��=%��>��D�AO�V��)���7���t�u��Z`=��@o:u�OW��*E�k�Ȟ><�7Y=�z7Ǐ��f>;�u�9@���V!�����r�r$s�7L
��)-��u�hY�I�{�P��Q���b!?�qz�;�(¿Hͪf�U/\��Bݵ�RQ��W��U����,8N�M�D���6�w+�T�}:-�NiV0t���8?�B����0B���Z�nt�{�x'����HaLN�]9���p����B��l���2@�ߏ@_��N3�S"���o��+^5=����"�6��zW�'@�c��N#�ע��,���	Vk�i7��E:��B(O��x�Z��)Q��V�@0*Nï$��.F:��59w�i��p�LS�\):��<FRt�n6�(�Ik��	�n��~�ra� 9A����PRB���=����G�P�ìV��H'��`��
ؙ>���c��^ 4{�|��aHؖ���3��7��FfM6�l��At�t�4���"[�Wp��]���yi��L��r���@ϖ����xޓ�η~�ȔV�Z���0�YQp3�#�7	���� ��T��jA����q=���I��3T.�?�Y�� ��'�Y�Q�A��=
�,��� � \F�L�Q�2���p"�n�>�� ��C�dϜQ�eF�j�2����m.[͖:vWwCGq�)��3h;���,_˷�M-���;Bk���	qi����ݰ0xZ��5/S9�6�K{n�c-Ee��}�捋:=G�<׳*�nfX�.����(���p�g��|���:C��H_�Ө��p޸�����]d��:���'c�o�M��J����h�f&G�_Q�-Wp#�b�⦪�4�e������	9arO)�5�c4���U��I��2�� 	\r\I�ӣV�u@[�G2Ot0�W��9G�S���j\�� �	[2C�,�?�`���D�?�˼��O/��u�ҿN��Ly�R>`�AM��DU-m��[̮�D`T��N�>P�+����B:��a+lL�-��~`7�g�W3�O��O��a�"3�|����P�⩒��?=԰̨DO{$d��4=!�_�
F~|��0aifI��`��5U㫾Z*w��י�宯٠�]����x�>
=Wwl/r!2���Z�߾����\�-��ھ�����A���u�Va��_�(M���R��??�l\y�:0Rj���y��0L*L���$`���:�M>���~2��]�P��zs���8�к@%�� v�fH_׵z��b���v��8ʻ����M}��5�8�~M��?�ZȾ�g�H��%��(7���|�[���|Wr'�ݎp�[�v��V@��^Mi��I~ϰ�=X�H<D����$G<^x~��pӬ�m����)�	�2�c�t����9�@>9xe�6&G$GT��&�U �H�h��2�~Z��Ck;T��/��	=�ij�]g���$�a�߭����^�e�y�Va�g�9%�L{�e/8�G��擐[�L	ף�iZj�v[Ǌ=��KTGс0� ���az���+�vSI|�?�e����ZŇ���?��w��.���7fG�&��0�&e��Td=*`,���Q�
��.����[�<��jE5�C6ā�</N�RȰ|�-y�x9V3���"���L��G�+��-��B��2\��~#΁A�ީ��2�!��g)�_#
q�o�E�Ma3I"������K!{�o���K5�<�iU�6�}Ohc�$(��s� D�q��W9�n�_
���BF\��H�!㐈.�1�S��mRdv â���_��/mmE8s�_,T��T5u���}?�6�����E�W�7�� �O��hu�}b���o2��޵#�	P�(�xq�~z�����>��5F� l�AQ`����y#��	ת#Lԡ���B�q4ļ�ٹ�e' GU�(RX�删�f�Q��5wKԭ1�A�Ŧr�!>�jj5W\� Ή�n�&�����m�	�in`!���I��?9Jn�Z��ƺ��G�I9���Ӗ�p�(��6�����ӷ���	m�*Q�G���߀��F��hzb�\���F�m��=m�P�;�㢹�慲�#Z����y���
��_t�FP`��o5��NK�E/�ܫB��A�*+�2V����:\���(�l.ɢI�~n��buJ^T�?��w�[����A�	@Ҩm�5��"��2�ɜL�� ���x��-�L�}��Q�+N�@����n◂�p\��5,�-	� ��r��D����L��"ҮHW�&��������;�|M�-�w���	���	|��7e�NL1��l?��i��B�A]���x���L��LW�
�I�#�Mc��%g��� ?�������%ɪr��0"�����6���$����f3��"�x�=�L&��Fy�6A=w���Bgz]��r��E��V}�'�er���r(�t��j� _�z��+���9��R"vK�qg�o�z	�Sh�ه?7 D5lOs�w 	J�8u�	�~�@RJCD��r��Q�=X��(엶*/ �Yl�R�7@B�I`i�F�H���^���NiW��H���'~�p����g�[{C�IW�0E�%l��#m}N�Y�<���S��<�wFDĸJ�A�J��}�Ǘ"?)�9?Ղ�c�U8���t�-���I	{��8!'�N� �ꊰ�{s�sG�ki�k�A�י=\��&%�ڸ���n�:����],c�ȭ>yV-���:���虎��n�#�H��9�2��P�Q�~uw?5���<�x8e���N@z����&N��*9�%���� �� <����G��w���s�qh+6�#�f򧘐_՝����+��Pw =�N��{�'�TT�jm1��]Zi|1�@�2������5w�x�pE@�M3]��H�!V��wŲ��a�`%��hc �:�㏠c{DO�R�,Ͼeu	��5��AJ��9�$��7��J��.'���-��v�o爁hLl�VWe�V�}vYc�xy���G�;d�4�!3��U �(_���q��]G˥�o ��u�6��!����Z��A�m�9�Ńʢ�XZ�Re��`�����N�&��0E���Q:Mj62�p(kM�/�������ɔ�M��o���S�AO�ӊ��C\�o�r�8]��	z��,�5Ts[�E���'��^��5�'���<��¡iL+$1�7沱��\��a��p��q�����VB�e!�V��&�q�Ñ[d)�����c�q��|��
����DF^1!H�-[N�hg|o�ٽ/������T�qB��Xmdt|h�^��K�4ᵽS���aL��R��x������q��}#>Z�Ĩ������c�e�l;��#$[��Xq���͌ �	���������r A��"K��W���#�����`�9���]��Z!�����M�c��S@�/�5S�����ᶚ�#^<�l��l���cXq�4��ZE���x��}	�P��T��o����v�'���(��w���v���=/\W;�%x/��@��i�+���Y�A����Vޭ&��肱z�����w�������-â��=[d`k��V,T��]�3�
��d-}��:��/��+ B˵�e)K잓��u�eM^�6m\��~���#:�,�B�ن��a��Ѵ�m"	���m��׵`�(q;��v�v� �_��r�:�dN7X�dv��J�W &��[@7�Zޘa�ej" �H=R�!�˒���/=G7��=@��P/�~M�����w��;�W���;���(�GT(c��q�CE�z
��F�{0?Z6\1F�BA�kw�:������q��Θ�:��[���ݲ��5�R��P����h5��&*�M<:y AHӣ$�-*�Q�c5!�f�c�<S���L&2*z��7�:��0�d�mI"��XX�n��xu�Q�p��*s��%����t��%�hMj?YXw�J̦]f�@���1���<������Za��-�G������9&���}���(ϗ+�-[ƹ�o���Z��8�46��׆ƨg��p��������$�̶=��ĺd����%��F�kʙ%}��:s���I��>��c��i�s�~�.�o?���`�6��9���{�w���+3�xl�:.��6i��	@�湊M���$礓S���E� i�o�6rM�G�nuϹw�/aZ��@*G"�����ؖ�N��W[��c�++fԇl�����|��5<*ԁBۙ�IH���-4 ՞ �g\���ߞ�F<�-\>U�u3z�N�3��S~ly�1���� i�X�����f�*�E0ԑD/aR��>A/ڜ���"=j/��+20|¯鵛ͻ"`����Zh|�Q��Bc�����=r����4�� �6E<��8{����?�X\ҳiW�s�3�,<lљ�Η��N0Y�����ۛ�kܭJ���$��X����>x��[�I��C�H-`���R�wWO��ď��%GY���vH3`�����ho�˷3j�]�6}]Y�!�Au���%���P��r��q7�@�!m¹D�b�uu֤q�S\�#/i�?���<s� [���O�6�B�������=Oju$rl��|��N�� <�c�D�Gô��r��G�r����*1�5��X�$�S!㬛��wN<Z�d�>�61����zvo�*���q�̖ ��_\�%=�
CDeSm:�2lĞ���=�Ѥ؟�˧x�A��ןG��Br���;D̯亵9,t��#Syދ��g�͛����7������/EjX8٪A�+�~���'�Vo(�r�C�	�\�;P[�f��_���H\"�r�����19,դ&,��	�M!�S���-c%�6k�����`�%��L�q��B�ʯ�`��E��Sx���"3�2�D��di�X%�%<v>Fi���&�o�����?�wz8O�����w���Ё,a�B�����~W�lc~��n)X�>��04��Qb��哶ny���c߸��v 򟐫(2xb"/��Jm�\R�+�o՞��W����jݴ��YQVB4��2�>������֚v�7$�'�~����~����OB-6P h��*&a{⍔L5K��¾�M�6?'�«+�ú8����p̄c�a_l�r��5��s8��5�vjz�1���?o�M�đk�i2h�ڴ�Q�F���y�5�v�@It���C�C�r$��&��Q� ���[(�j��a�mGO��X9���l�tI���t�X��tR,���8�v}q�9J�tyL�YY`f�����c�|V9����܂���M��qߥ�g���\b=5�����27&�f�Τ�W�eh�U���������M��cʇp��
��Z�ݷ��ʵ��R6��0U/�_TKv@EdL^��B4L�)(*��*�!T�ڽ\>����g�r{�zx��ߧ�'����E�8x���S�e]A@��(6�Q� ���C��hA�5���ѹ_8F���DW�1��(	2x�LB
u׼�8��7M9���������a?����μ�҂&�X���؏�嶋�XCZ^��.��F׳�R���(�H��o9l)y�4�q�+R+��FA^uڝ �k鳁4	�~&��P( ��!�bb�����' ������(8a"�B��WB�󛅖��aZ^�.}��kY�
b�8�n�o{���8� n+�lo�ՕT�<:����=[U44�z��XFC�ך�X�?�?0�Ծ{�A b܆!p%�N\K��Ağ�Y���N�Q�O����3'���nI�C�O�c��}�X�;:�ѧ6���wg̑���@/�(�{>=���y2�$�2'��Bw��o�7K%�f��Uߕ��3�P-n,��jW+,uC ��5�`2F�m?�GK.ְ�b�d1I^�p�O��7�@�>'h�ϔWO!T~�#+Z~��}ģ��G̰�>¿��dq�껌Z~_�����b�İ�S=@~w�����:�������'�єg��2�)��B��m��`3����]]@�E�����B�a�bs{l�ز3a"Y;]y�(ec���xZ@�)�$	v�%�ױ1s��y`� g,l��?��Tg��z	a���:�3f��2�YE�jǰ�ќދ�Ađc�5���*�]\Ҝ�ٻ���i_�=�+{�7-� y���*9�{�h��3�� �ʀ�"�|(�[e3��|�ﭰ�b�n��?5�ov��%�OG��\��	�`/ �r���o<���@t�E�X5zޒ�t5
�ً
�$�XIZg$Cƍ�Dv��u;��c�<ARK(��FS�
�┉2���7��6�� �9}�h���\� ��_�ot��8^JV6Sv%$DG�D�|���6y$�W#��"���V)N!G���5C�>��۝@R�^h0r��h�X<�S�C�U~p��u��sB	S�C�ֽ������&xѢ*����I���y)`ѐ[���x�lh�L�o��
��lA����29�V�@��)$��3�x�1P!5��+�j�����97hK.�C��M_)/��|��ū"'�F��Z��#���?����:�������.mD�"q���V7
�K=��<Z4��(i��;dM���KQM�x��%ǜ���~����a:Л0|�Cq���>��%��e���C&��,�{q]�I)�m�S�6���@t��Nތ ��
w�a(�\D��_������M��]��b���/���eVIܶ��	�)�Pm��:��M"�û�\�t����3�m��"6�^�l�L�F�Т���q�������c���R}�X&G঑�ȍ���>W�K��ƙq��'��Ϣ��l⨣I�~
^�thmtM}���6i-!�T9��<�{�۟]�+ �<�|��
͋��N�3�FBß��c�?c�;���θH�	w��?�O�!h.�F�<�*�b����ґO�{&^=/��h����f_�ҢL�1��C�iQ+���:��U�	W�BVc*��(��ߋ�៥�s�}�6���t����V"�XnB�����Z�S#�����8f���c@6�a=��֭���5	 YqYZ���4]Le��(��/|f>-���kt������M�v7[���Y��i(v�lɚ��GB���L0%8�2Eڱ��j[�:�~*`n"���#���d�$y��E,�����g�*�{ �aL`t�9@T0�9�Q��g�»$�<�A�Z�.��t��d��ޯ��415�V�R�ܫ=Tى�/�����+�+�C�{��2�ĕ�����i�i��@�'��<�<��p,��3�T:u�,?�H���ȺUㇷKH����x�9�������i���ϱY+k��wt��8K�wCn��}i &,���1�g9`��Y����K1�s�D�w4\� E��Y�%�x�Uc�Z���tG�X���ex�2�AI��v���T��8b��+:=c�u��.=�j,0��M�LF/�`x��"?���b��^�B����B������B��֔si�������i�eR���Vӊ=�4o�O�_�;IJ�0A#m�ܣ,�U��<�j���PLݙL��y%�i��n�4�W��0�N��~,�G�x���7��I�ۭ��� 0y@�{�N��#�$e�j���́�Q:t᫑zp��(�o0 ���M�j7Fo2�	��M+�`ȯq����lM�����H�w���Ǣ${O���^�R�^�&a�1�:e~ �����eY"u��Z2��DT{ ٞ��-�W�p1bW�z�{����aJ@I��D�=ȰV��wfN@�_�7�������N\E#��>���g�