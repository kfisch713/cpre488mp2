XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|%|���Ѩ��a�L�\�A`WԄ>4$�2�qVyp��J�D�� ��3�g���g7�R���$O	�Y����yM45,��ֲ������M��@\��؂��F�$�)��$,.�_q�+(�L��3j���7KwY�[�{n�g��P�Ӥ
vQ;�)"�z��"g���eļs�:BҕBk/+3:�?@G�\�G�,nj}�nEG �WÌU\�T���|��|[�g��N,`����.̪5>�(�-<�P˃�t�b,���P	��uv�N珮����4����$e�\��`�q�c�ɵ�o���GCch��<oԟv�zK�\$7�>y�����K�4�݅��DOւ6����M�7 �P;��.~�H� yB.�*��J��n%���p��&����h%0g�v8�q���}��E$U>�$��O~ǥ��E�l��!�c"��v��#���W�)�)ƯC���ĦBQQ�0�E�&IXF/j����҉C׫�_�?T�&���2$?����wg�2�y���߫�i�Q���x �.��x�A�J?p�X�T��[h���]��~]w8���ȉ-]�	3����,�qĔ�c�=�D;#
L����F�3�S+�c��&zũ=Nj����� 0�9Wv֢'2�K�OS*�Z]Ӝ�q��3!2��������I���7�1g��ޛS�w]9�~nGu�D4��*kߡk�ct���R �[�.=�;������ʺ��(#�ѐnX=��*v�����nU�B�ɑ�f�HpXlxVHYEB    241a     ad0� �3�߭�T��}H�{|#�Т�9"��VV��xOVK�x�d�q-�#�3�m� d����
\�:]d��j�n��v��`��~��*m�'o2�s��֋s�y���P%�K�d�=�$p�iJ���_����`�z@8�ɹ�RNd�Hº� zTƄ1��ɢ z��,]�n\m��oA� 7��W�jmT9pt���%M���ѱ���{wZ�1�u+��Õ0u�S�S��q�0�0ڻS��!<&�
����4o�B.��)׼դ��0�����$ǔ&�['ݛ�����b���p"b;��V�:X
��v�����}��.](��*}	oo�m~{���)Eqi0(�%f����yα(�� ̥<�$i[�����&*sn�6H������"���P��~���>��-�mW��S;���1ͪ2Z�V�"���@*�>Ix����:�*Q� 3t���н±&�9Gt���r�L�Ћ�Q�Yk���Oc��
0!�k�1�F���w졼�hm)e*˖����qa����2��Pk���S�mk ��������Z���ןߘ�S�C����(>U�̰Ծ�nL�8#]QO��ul�Ɋ��p�_LF��>��S[ ]��Y���<ws�J�C�w�1	�W.���=�l���\����l�mZ���^~�fR���b���eİ=FR�7Ɣ`�0�lw�!_�����Y�+�zK����[�v2�yv���SU��ajP�@I��ݯ�n2�<���3�$��6Xi��eM�8������H��_X)��XL
c8t=N	���� �=f��&(<��(t�M�<m>h^�'��3+}AC�!5.UHKت���K�bt�r��l+�b���Ar��Rt=r��g����%�h2�
��\ �.-c������n,��r�C�c@�*D�\�*W՞�$�;:����fה�m����}2����ڷ+~��p�5��;��[���!$����p*�C^k��k˭n�_�9�z�Q���_�!E�_&�j�e
��nоpr��L�M���\Z������@I�ǳ�<<8)H0�R��a�H#�&=䟷���
�j���K�L��]���:��+*��d;#!��`B���f��Z�s�3�* ����+����!�`_���U6��mu����4޴�����zo�E>_L��IGӳ7��O�w�N'ͩ$��
�~$b=�@
t�bդŢ�ĉ�G�Gl��)=����|Bo��d�	I<�珛�M,D�e��	)��ཽC2����ϕ*pK^Ӈ9hy2j`�T.�²���s�z���s���)UJ����Y�g_ec`A�y���2I� ��(���|��5��1��΋.��4lgO�z����b�\���3A6���0�{)�~MQA	�Dmۺ@�=�uVߏڧ%;�������y��2ݫ��� �`�sŗe->��<�XR�'o�w�HK߸!��t��x�\~	�e��6��L+.��KAgBSf|ȱ(=�E�ğ�)UW�g�{� $iI����A��!�S��e���3�g�	ъ^��ߴ���۔�-K� P2��	��:��B��Lg�D%55&�͟$]~;�0�6D��h�T8��jf�]߮��#���o@Kyp<*��U;v��t_l)�J'��\�� �Y����W�%�ZI�)p���P|�3���Nrx?�AT�V\�?�I��E�G��ϭ#�)>�h��z?���+�����.���?˅�k�V-�F��sܢ?��34~��h	3�����lA�ml��w��:աP_\S��}����Aq]p�E�8��-��4G��i�P�ܯ������+�,���6���φǻkj���X�ȷ��lң+�>V$cQ�=؛,�f�1S�'��J)�OZ�1��&�X�C|�u�]m-�m�o�z}�8�a��s���ѥ`XL<���}c�Î���x9u|p�a���GA^JFt��D�H�Ю&L��#�S���;���ӳ3C(%lͣ/�/��X�{U<��p97�D�R�,Lପlw������$r9a&�>����I�������g/�s��W�=�<m"��T�
ͻ�*�lM�r~qj�d�N�-`�b
�#e�4fO-��Q��z8����0@=U��A��m��S��[2����4$�!_4�����q�Lx�%�Q�5@�g�l]�xwr��w�K�����]]�����[�C~q�3�ﳵv�]B�+����v�*�h�W(�ړ�z��O���m�m�z�>lP+	����qߑa̎�K� ��"�b�=i"�D�YQe���z����F��q*�t�>�n���'I!��0�5,|+Dt�+��<�̸����q�fS��ف.��d+�X���$Smϓ�̃7�>��21.�=� v�����CYToU31��FifG��\����gtE�҂I>���
G�L�4W���q�wͫ��ΥV�A}Q�gR�� W��k��,Lt��RjcF��T�adLrp�dķ����钅o�����Q�s:Ue7���ś�>r��֨|�hj�3y�U�����*~'��.����KC2����nSL` b��?��HW�������G��Y�];�����Kw:�B�d����!H[�	�p�k*��we����&�Y��G�֐&UÕA������Xy�e��0�ܸ>pT�����A�g��O�c�>!Ͻ����V�X=fe�R�