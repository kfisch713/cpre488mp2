XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����hi��(^�;�����W{sVj�N l�8��<��$#�oqP�9�ϊ��Tx��{oٲ��?�ezZ,�;s����u~"V�W�I��hg��摚x2{��4�
�������o�Dj�mC�`�"��Ƚ�pZґ�>����R{e����k 
s<�)�[<�,��{-~_�-^���D��v�uO���;d]��Z��*����ٿ�6vw�]�/��W7�q��@aH�=|�,�,3�!���� ��X\�q�������RB�l8kf���b�u���� K���&��7K$��2N�	Kc�_�8eΗ���R�i�y!!zZ��M����#�]YI������� ��ǭ��7��E�xSt����L�,���݂1��Vb�e��-"Y��O[�?o�bi�XH�^���%�j�\ϻ%���3�?������E6��	ǧK�NM�Ag~ 0!!z�ɕ*���)�I����V��@�� z���]A�'��e�b_U~|�e��}�y�;�P�W�[W��ӥã�C�#	�3-UɿB7~ӑ�UQ��W���.���?f信(ۙ�K�ᰄ��
��D��|���~����l�V�z���l����{E��,�=�n�1O܇�����7[C�L);�r�����a��C��V��S
�7b��ڸ�̥�"����2u^�"�������Bg�)}�ΠT���|��B���(�4���7�imO�7����u��@�����Cv�=�>�HXlxVHYEB    374e     ea0��(��o�'T��/)�:C��8{�~mk��{��	te�џ�vԬj��"���f�}�|pч��%��'5��3�� ;\>�`H�����w�)7��[%�w~�F*0�UF�'@'X�C4,w[�9@A�XF�u�7 �{�
V�G�w��o��W-s���Xe'�Y��t#N��0�Ky�l�\������$�9�|E���O#a�ҫ`%���*U�_Y���Qƕ�~ڸ�b��JDҊm�4K��2�G�z��� ��z<~�Gi"������"3���enM�����>�����6u��	��4Q�^�@���Lq�<dn�x�Mp����\lw;9�HzBk.g,1^�f�FhY�b
�:���Ri"�H[��uXņ�Q%	'2��S�}�R[4ӌL��DQ��ո�؋{�Y�L�$ȿ����g_�9��V�Hژ.�D,;�:��T����ʇ���s��R��/�<4���p(�Y�v1D�Dw�	����D*|Mt��0i��|�/�ָ5���$:���D�.�A(�W�i��	]�G���v�˧���c��R�z:�H!>A����l�e���R)?�7�6�Ր�
���b�����TKb�&���h0�W;:�A�ۚO��D����]��I;Y�@��*|�ߨW"�<�צB8u?�x��)O�Q�OK+Ϥ �ȇ�F�����4�CK}����8c"�����әC�ǿ3Ⱥ�%��9Ť�S~Ȱ��������Ε��xJ�4��$^|O���¬2��9��5�cB���q&tЯ�2gS/54?����R>�u���E[6�,\Wcg!�4�(��ݫn�jT ]�W����8�a,|�y�奁F��MD�ǟ����%��|����T��}���w���*�3h�e%d&u�9C��سM��Cȃ&��ϭ���X=R�' ���i�� ����\9��:F\��%��8���U:���[�o�t�K�@)�
�A��!�W���L���V޲j�;�����4q�$OgxDH�m��5���� g�"�ݱ&D̳륇�QJ��"�d���� ��Ziy�X��x�a�n�-�*�س��?�R�g.Y(�T�<��͠�>A�2���Ǜy��Wƌ���t��dg����3U�Q,�Bu��W"}��Xo�2h1D܆�
Cum  f�<��$-���.�
�rˎo2�n�~�ݷ���|l!�2��I�*7P g�ѫ|Tp#���L�h2KH�=�N�n�G������y�מ�n���`QQ;G��T�&F�!�j��3�U	CǚNH��"�v��Ԑ�Q��5� �I���Ɯ�f��H���PKV�p�n�p2�������7�D��9�|��A�<��huӭ���%�[X�i�u�JV���'�Wjn.��t7Z�v�S9�t�SF��I;J��EJ�'�v?�)>R��5nF;�W�>yf�'��*���M�":��$�YSXC_1���PK\<���|	M�x�<_���	_��`��^IA!�u1	]��0&��&]n��ͯ�=Y �yZ�l�qW__��h��~������?�-3���vc3y�hS<�vr;�b�AW!t�{|4�@b)��e+�괛��iC��r	Q�q���P������H�)۲pď|U�"=kE�9E ��ˑ��C���QC��RB]R����{�I<N��C��M0j'b)~��I�㢐HrqRעy'ʊ��P�M�f���RUB��=��2��@�:v�,E����.�M�6�4&�b�Mu��Ś� 3��� �j,޵�n�?ϋ~j(�r�T�������:}]��m-U�H%�L�+�����:��/��8Z���C�@�+=�F��//m�U����b�3H-�H-q4�n�_�Vc:Buܟ�� ��rx���0n�"�W/HS��@(H��:F�wcgr+�'���\�����JZ�x2�%��ZЂo�,�O�>�T�X$-,�,�}2(�������kˣ�9��l������ly��ݫ��4o���j����R�_&�N��*����u���k�K�,�����<7�� L֠�az�C���Cf�V�tC
�3�4Ѣ�W� ���̡�����@bˁ4/�V��3i�\ ��L��Ь ���k��йi����Όz��l��q���:�5�,��τqmbf��~�׊�c1e�������{�$S�ѫ���9�,R���q�$ ��t�+��CjH�8�7�\�qhEV�)�Y�ɋؚ�E�ؕ����\'�G�Ѕa;��~Mqο�>a�H�IQ�z�jߙ獃^��T��{Ԛ"���HjiWZ�Q��UX�OȨΜ����i����h���u/��mm�.8J?��oa��>�����5K	5ȴG� �ir��������"�!�4��p��ÿ��er���z+��w]A�6}��?vؘ����7���Ps� ]ߌ�P�������n� �,�4��*�q�]��?!�3����x��}Ǯ	� Q�B<o�"^M���P�Փ�,��`�1��ѓU�`��v>ycT��M|W�&��K���f���ӯ�V��E/@ ʕP�ӿ�����g�v}>���Crd9���W@���ô,�P������^�=�Z�V�[���	w"j孢I�hY �|���e149!���<�P�KFr���ʗ�*_��\�a1����yf�zE�����
d�ɠ`��O=��޽�!��m̴��"[4>gt�S�ʋZ"���J Z�`�q�uq��*�Rx����`�o����6��x_+�M� w�A���ˇk���N�m/G�hq�(�+f*�qMYW֍_���� ��H�^���mS�v�K�M�%&�2��P/���|+� m��?퓭��./�Y=���7�bXv�]���[~����Y�_�r��ܢ����A�5��b�p��o��'�9;}h��e��W���0�+��<�.��04K�=he�5Ņ!t9ol�e���1��Q�N7>UY���"B:�r�������v�N'L���~z!m֙��=��n��>$�W�݁�4��x{�_#U`B;���b�}R�v��n��m�-e}x��y�k�aҤ���!�V �A��G�;�
�y���fpW�*v�]u�(��/������,�|(ی/���'�F�ORlZ��gm�4�,��n�s���Lrǭ�t>w�s�0)��0��F����;�+K�:����F�ο�r��3G["FYF�q!�B>�²���K�I�C�����U��������z���$���ijZ�:����{�-+�A,@��P���HW�g����F�D@E?���6/L���mO����g"������&��k��.��
��0��}38C�`�6��n����=�P�Z�4��"�V�.����#!f�V5����yu��U+QY���`����Ld'��'��Z�?���8���m�-d�o߃GZ���{Ӧ����W��*M�W���2�� ��90E����D�����8�L��>�r�z�_'�x�Paq����ܰm��
ϑ6j��c�F�|���1f�j.���	G�,��+�B� aAؼ
l�N�	C�-JEq�y��P"%��&r�*�~lErlAP<�8���^{��cV�}+<���1�ؚ��jJ�65��e/ms�Í����d�����!�Fs.h!�"-#