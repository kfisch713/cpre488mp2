XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����h��?�3���cZ�H��?�Ą+$�4��e����0W�:��?��Yrc9��ʮ� ��Zi9��1�7�[��a$��(vÂ�0~���-'|MN���yK��
��)mUnbZ���C�ʗ�r�ak{�k��@
���ޅz���M��O؆�nM�懹I&��j�����U}�W(N����6�t.��;�yf���<7�����y/����_������𞌆�/��:<�I�E'��Ԓg�CJ[	������d
�����%�:{���Q/V-�� ����a\ndE6Hv���1$��iy���UvJx^���<qN�|��n������y5��_��c�����s�}��Q`_����9���"��KA�fv�˳�]|�ݿ%���ڳM�cڙ�z�&0���������U~gi��'z�9&]�M�S��b�� ���3	=JO 9�5�ꃃL@��U���ˬ��W�q/�'��-\[����ω2g��t:P����e��������N�����<t�,'^��"��-�p�iX����U9�ah���+��ޤ���E@���'�A���T�Ax��u�ԩ?Htb�}�ŕ��	��Ϧx����y��O94�K^���w������(v���0��qr6�L�H��h=�Zo���vޝ�1�ǟ(q��#�Y���"�k�j�E/�A�+���ju4�_��E6�?���
�]��g�EJQ�1z�:k�f�b�X6~F��m��8B��O�4�7Թ��LXlxVHYEB    1853     810�͕y<aw)J���|Iԯ��K�l4�@���!��a��������5X�kl�t�żQesf���C
{���>R�.:z��j��s��1�B����� Q>o�*�R-U4,�5z>Qy�F�.�c,��<�s&xi���;ڱ�7�-a�x�������8 ] ��h�U�uMi�س*���g~������*wTNE�	��g-�\I9j�ٌ>d��9P��G�;*��q|^����t����"�����(;�_��M�B�\#Iޥ�� �]�z���p~~�@�%������n	>�q]��o�[F%���Bq^Sd�V�'�_���L��F�M��9�#L�!\��C@��� cK�}O_�i�t�2~ꗟݒ"��5���g��%p[��o��j�7i�;��Ya��� ��p���hE�����x���/L���SS��3.d�z�����`r�v2h�����>����m@F��=���p%1J�m�:e^r�O��|��p�I��A���`�n.�]@9�@�:�+Զ�����B�������	`�ŌRg��/U&�. F�������24�����u[�s�;\]�5��$%O(|��	E��{X61a_)!K��DA���b���}K됕uL��<�Ӊ��qH��@�� +۝#+��*�X;��]�zk-���q��!��ڨ���3&+�g0���׋8s̻�ŷ9Փ=�x���(�ĐjT�tW�I�M�{~r}�V�Ki笰s�E�H�Ê��1�#6ȶ���Qڌ��s�@/���y$��sW����:���+2]L#�SƮK�x ���'r��G�����W�Ov��p6p��f��s�+��-�ݍ��\Nt�T:���-�v��CK��, *�ҋ$���|o�G��d���ɽ����abi��qZ?��&����T���dj^����@k=Ss��BFcK�C�j�Zr���K��-�`���Eܚ]�3L�l ؅q��@������� Bg�`)=�*Ӭ�튓�0D�j�ԗO0TO�JU2zG'$�Sȶڐ�eMp�����k,,�V�XG\�_��������Y#'��a�(��6-�5b����F������J*�Ғ��a�[G{�(�#(�J{��	�~�/-��7�lp��wnu$l>;
6Zut�4θ
�f�2�pX����Ӝ�[�f@rv]i����7�x�,�n�a#.�x�h����ĭwg�P˗:��u�X�v}�荥{Ų��z��=�O!c]=��ִ��ߨ�?.��8Nϳ�Vi_o�Y�\J$�+����{d��*����R���)����(o�r Y�q��+��1X[?��{��L�Q���I����*��u���=���;@����E�>�����oJ��x�WP���+��¤���
/���Fѣ3�[z_���Z�l�!	:�Y4�f26��h���V��K
�E����4���v��`v�G�o�-o��Z�M��Pww��4��A7�9�?��fU
8-UZâ������+Ӭ^�g��>j������/r*�o �m�
_��G�Ѷ�`�\�����n2����V�� N��u�
�I�Q/�5�&A��#S���cB���e��C7,(�� ~k¹�|�ڼ�5��y�^ׇ��1׷ce�&Ң���ֶ앾P��@%�-�%cM����n��u�!�T�	���~2�2X>#��������)���A��UE!�l����&���G�wD��L��aD���揃K�x(#����3�U�a��2)>�HQ��w2��8:��7�H����b��/�c�~�uĮ�a�Y�Z+��P�TA��?�F��Z������Vn��V@ ��_~���{O��P	�����p��͛؍�ųpZ�!��ޓy 9��ϒS*!l>5��&Byw�������T�<��{��6��W��]E�m�ͭp@��)�tq�E�.���6�����N�r��éZ�����ՒЛm}�����m 4&�ϫ,�P�zC��Ղ�d��E�'��(fFx9!y(��