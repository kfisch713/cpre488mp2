XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������{.ku��X[��<��X�0�y_��*
l��\�*2�I���TZ���y�S�@�
k������G߁G��{x�}"�Dvz�	EB6��Ôr�3홺�4�r�_�%{;l@ǂ�4y�U�^���	I�3�F�@���O���d�`z�IAB�;=�B a@�U�-~�܀�ƨ�6��� �ʈy��Ig5��$�$�v�� L+G"�	4�(S�iB�D��/1(��f�eDB�B�����@�r��HJ�U�lѻ~���5���*��?՗�@+&I@޹�K�C��d��1����Q���B鵳k~r�;�ù��(�����9ȆE��W��k��P��Akq�g%%f>v�ϠTjeAKC-�ή�a�4�&��F�-#.��8n���4��]%ˣޏj��uǾ���:�qrT�ksEV�Y'�\ƫ�� ��X<{7�찀'�����K}P�}�8�w�B``�w�#l�9+��I��W��)�'~ ����[��B́X[}�Y��m��+�í��,@+$��Ηݖ�%̯.ݲ�g���~=+R����)�ݛSF�qJhg3g� �I�S��f ��N���t
��R�*�b�$�Päte�*�ֻ�ᴑ`s�d��2�~�~�|<O�V�G�r�$)�����Ex]
�8�\`-�m�uC�w�u�l�1 ЛV`I���Q���K����jq`p�����Eզ��דŚ�W���%�(��:�V�XlxVHYEB    dd8f    2160>��A��K�!�(8�9k�K��>�H��S:,���e�R8x���7�D�X���qpqJ���K8�������Z���y�k��p�Y�}�&���3N��}
�@O�budk���q��*a�*qjHd��fT0<h	e�8=�G�b!�d\�g��U$�ښG�>9G^���,-;��1E���-G���@jQ95�����"|�(�6ǚ��#��w����T��o!sCS�_F
Iܥ��t?��y�Q�"=���i�,Kj8�Fa����T��$9�q�@*����$r{���P�qY���]>Ңe�����B��]���`{c����5���T~<�c-�*�{�3r�~U��'�F�K���e^:��ѣs�����wb�l(��n�8��O��ז�X �+���g�p0�'�V����mX#��Z�o��J�n���A�8���|ɦ���h�wu�G�+IO+K2�+��Q���2IID�]��}�Y���Re=��!W�= ��yN� ���S�W\cQk#Ē,s���f�$��?�B�����X;�(���Џ�I#�.YR���^m*H�>AV�.3��%�;R��B�W묊5<�9&|�\�/|�+�޹�}��E��y��)������o�z'�Mh��а�d���Kj�!B`�gk�bx��2.���"ck�]�����N�=P�ʩ;`���A�##���n%+~X��.��+�_��Ӕ��)��5*� l|��>��l('�j��[��˄8���5�w������tfm�J4I���al#�8��hx�iY-ER��N��@ ��"T!�9�(){�k���Yc���K'�MV��is�d�A��p7WWCt4g{HdA~���'f1�2�W�J�żB������c�R�"!ÂQ��2�umiW����NfEm��f��Jb�$0�PQrz��&k�}���O4�Z�σO0"��c�ؘA�4��7v.�і�3�8�p)�Ҫh�-Yx����=Kf�Thay�=���S�8���"L�ڊfL��k0���W��o���v͝q2q;#��m�]U3��)f{@=��c��,��	$��/g�DJ����&��%/��.�<�W�-62�jgPMX���/�M�.���3�}wE�����������ߩ>![Z����,�����ϸB��4�n���_��zT
���>�<�v*��s��އ^��{����qML$��Tr��4��b��Q	�TpY�$o�WpnY��2i�k=E������_�cP�Ԫ�;��d �� �s,��XC��l������Ȓ �����d�"��n�C���/���;(7���.�+Qꌞ�o��a u�i��Q1�Il���:����� �מ�˪��o�6����oS�1��_������D-�ɯ�7�����,�ѭ7J9/�2��=����.��Q;�j��ܝ�j�vk=U7}S�*Slxh,�l������3�!��
@�Z���E��3�?-K��x�k���t�O�>̼�u�L�k5X����a�XW��Bv�jZ;�Qet�b7ŇO�`h@���r���F1�R�3䇚����\����&40�4ڸ^�����7@�	}�I�!3i%���k�8�h!�KJ:��m�2�]%����{�_�4�}�̯�K٘�v����2����5���^��Y�hҶ�c564/.~����u��ՠ���ҝ���*����n�����%%�,�<�a��1Fh������BI(xao`�d���^��} }C\�1�۪i| �k<��I�*�������O�m流B.�g��������Z\��hk+Cb|����I.3ѫ�����w=)l����Ϸ�vW($A϶#�s�a/�g����RX���W��g-B�	���v��������9�Y�T���L��'(��mk���?
�,�8<x%ƒ�ix�Р�%��ݨ�>;��M�C+��w�l��(���I"JPsu�BF2i5$�FY!���,�����B�*7?�����;�Q0�AJ@ �,�k�i�+����F誇A6ڻv����l�пdE�d�����~�L,�#����/��
�{^��� �,f���,g������LD�(y��u���oH�D�ü�o\ ��h�bJv�L(š��ٚ�N/~��S���<��I��t�S���D�8vH�g�Ʀ����xIP���X�T@�j[��mnXH�ڟ�)�l�B?i��A8�8K�W͈҇v�
�k���n��op~��k���55�b�vt=��ޜv���dY������)��y<l�Vz�O�Տ��m��8�s6��q&7�OFV��6l���K�������!"��v�=�P�L)2�(y5�>Az`�Foq�`	H:]���EX`���'"���T�����S�̈́T��'�1l�G�T�؛����JYd�w�9=�-��=��m+>�����C�� ���]����x���ј���Lf^��ӓ0�1c���eX�/,�OwIp�gIt����M��o�"���U3��/�ՙ��Ձ�v�^r$cYIs~_�Qj�v+�j����P��O���!���:AC�]�ѧ�lp��b����n5����D?�ZByͪ|��-�<Uyu�nn!|�?���飶�c��F����yx�z}<���|M�!��yi+�������6H�������n�K�.(���u|�1��W���f�7�E<q��6����A��������i��hjh㝂)�t�ޗ9�$�<ĂE����z�gDF�Pv���G��l%ԏ�[�I�=#�����T���k���ga4]��Y�DI��e	X�8="�>�� ~�6��T�8l55�c���}͇����nmA�1٬�vsf�E�\�ͬX*�hrT8~ʻ񧹲���$��x瓲�E대02���Aڐ��(K�>�w�_n��{o�o�L�� !�Sb�'��.~��i-��b쾛�aQ�S�4F�1LȹC4o�PL��i[�U���C��{��J����i���mRnOX!�8w�u{E�3T�����rӸ��S!�S�Dl�'O�3���6=H��0�}m�y-0UY�'����}��3�%�^�%jۅp��=T1t=T�Efm2�1���R�0h\�ИxM�3z�٬�Ȳ*���س�gՃn�����z��ϊ�0�G�ك���;U=4�Y#Y!��4g&@����Q��bD�&B2҄���(��H�!�l��\�\���$��s���}+���$.�Ȏs��_�9at�="{a7�r��4p8�Ld�aT(jk:@P0�����<T�����E�V���B�������������y�p��2�	���rSp�ԋ��h|&���I3vs��S���w%I�""�
�a��4B ]e@�`x]�^�����d���F[�J|�aī�o:P~ަ-��K{'����1]��\�����#��B]$417bĩ0�f�/S G�Xs_����F\=�l�;!�M�`{)��-�t��(ݏ�r���0T�J~qi��o_IgP�pJ����������;X�uׄ��x�\ѥ��ok��3�< ��Zk�/P�� %JW��ʏ]��?�o�6k�9K{�Un��h��8A��IM�.v9^
+1�K*?�;�h�c.3��}��^3��/����(��W���{���4�3������������5�Lf�*�r[��}��;��2�P�t�a녖�-+φs1�L���<���݊���$�Qo5R��|e�@�˲�
*+�.��	=��kA۟z��`oW$���N��#���tÌ�N�)Τt�,��zJ5>i�L�Ǿ)l�Q4�T���Z֠9{����HC���4�{F+7L	���?&v�a7�,��P�pi촰��ۿ=�c��.1Z}(�5YY�P������sR����l)����|X���]
H�U!��"8TB����s&�i/&��g�#SVIrc��՗[���L��;���#��H�]B���lYqZQ�=�g����ǘ��=�=,N�a���]��u���5/S����n���	�9g�)\\�!�Q�Y�r=��t#��&cL�T?%$"�	�_�ޡW�W�z�=��<!�K#%��"�D���1AL!8 \�r�ˠԸ�ܡ>�P�dO�z2���������~uL��:kF�Q�(�������p�m��k�2���:�o����RI�`��k�a���qK��+�D��ޝcT�8+�_�0<�,�Nv=@�i�t桳�猕����_�x�1���%`�ZiƸC�<4wq�`3�լ�p]��B��&�}c���_ŀţL�������;���4E�Vq���HA�z5Vu]��:�Q4(�\şM4�4�0���xy��JZ�z+�ܗ��Wc�ᝈ�lE9s�j��җ�й�ɴ9�9Us1��+3כqK����o��b�bS��7�~	�Va�[�,c����-����RL���!~k!6d�����N>���21���A�/����Q�K ��<���F;��N���F��"(�$��a�(!G���qI؊�
U�B�O�l\[��n�gC���,������/��r��k�i �v̟mu��E�C�����W-����-�o'߱-@���5���,�6��/`��r�++z�'!P���ne��x�Jvw�Jq�[g�v�S@����*p�;"S�a��\D`�Pfn�r�����- &a`A
�����[���#����-�����j�]�pԓ�&{��̅Zӆ�|~b�"��~�;<1������~U�¦�M��̠W�7�r�E�������б�47�Q	hb?%u���*M��EA�Q'$�`mE�b�ةѱ�d�=����s޸���# �:��w*��KEʪ�bdv�f��0�ss��s�v�q!�f<lַh�����Y��A���\w������s�W�;�.��"�
�7m�z����E��Q
?�f���>q.$�b��A���9ё��6%��h�'%(�Tjf}����h����Пr��"�]�/I�8fbO���h�q�*9�t\y?��u�t:\���e�*�J��'�"w�AQd�i�6���J��?M{Ӡ���:�",�����bz6���'2��,V��Sn�BH�gS�b=�Rמi!��������f�a������Ko��.�a�ֲ�t	pz��D{�-��(׽G�����2\"�.�H�ڑJ��="d.sa.��m$j"0�8.�YUI8����8@4�>�|�gm�����i8�8��	{�4)m��f3��� 乍 �ľ�͹T<��əS�⺄��7�Du$"��d����	'�<Z����W�*EY^m�p�*�(���,F�I֏#\�� T�f����l�`:X�����.'��������ދ��Ngc�-�����lxFN�1��m�����h�0�R,&]a�Ɍ.��e&�G�Z&���\a��<>�q���F���b���uo;`��^��h�
r��R��x��gP�Jx��j�n7 `����g�֮���T�~�C�e�1wKOm2�� A4�'$-��gl����@�@�锨q~~,T��{f���+,��$��>Ew��V����7y���5+�B$�Ƭ��5�šӌ�Z�GoC-E%�L9v.i�LJ������0�[����dލ����Kry��}!�|�0E1����T��7�$_^$��Y�m���}�ǫ�Kl�m��R���ϸ<_��J>P�є���`����C�D��5lp��ai�	�H1����ʪó�U��,�B��֕�Au��&��;�L0����o�OJ��U�[��hmn�㘀a�"Fa�k���UtCl����׏�[����=�v���V�E�pCMn��
Y�s��+~��Xt*�:!��\G�`��d`*j.@�]��Y�&͔f�[=��W��"�Pj��ٰ�;/"{����$��N1���12>����LH�������>:�i����
�Ƃ�&�K�XB�<�;�x���ʌ$�鈯g��0N�W_{m���ВH�s�j4��΢�ꔒ�K�Txg��yi6�VE�%�u��=}2�gRұ/��l��\�b��QI6#K;^�~D�Y���u��8�h��Uڞ}�r_x:}�dD>>J�+�S�A�3�b����D������
��j��N�"G�6�^��B�uh6�rg��¨g��k˼��ת��C�6м �MC)mC�I�s¦x2����5���Q0������}��y�8�����̾Hu/������"�˵��{rE�K��ӽ��%{�_�þ�irMղ��[̽pV?�����E�&V
���`�e�G�����zg�r�y6�ѸU厭.����+��s�*뺈��G��.p��� I}��
�λ_�A�2��tr�~�$�:��=QQ~��C40#�2�
n;�蠸L'� (�T����/�ԙ*M�L��"9���+��.D.!�E�L8�xtd��b�F~�ubmH����N��kX�6��s�J��l<)����������kb-{�������a�O��ӳf��w�c��Fy�`+RK����D�|'I�g'D�_�6�h�mS������X�*H�ղD���Wx���M ��3����RIPW��o?��D���$�w���]V:$4��г���;՝j��ራR$�5���H�{�5��p����ѣ�G�������N�(�4�
{��~��&�*�Y%�/��m�	ʼFY�d��씛jTp���$q��WH�AhPDΎ���i�'3C���]�a;�Đ�j�xw�#��t�S�C����/^6�r���'X=�i*�,�&�{��ĸ���aV��-���l��F�y"; kU�է����iJ(��K"��K��Q(i��=ZMe]�OYs"tT�`�pkE�[Į9��>�s�7��+�W���o@,菾������}H��S��#\	�e(��l�z�Ř5�P<J~�Տ#�Ď���Ó��E�/��yM����'r��bO"@�ގ��J����t��% S�w��_r��ڱ��m�2&t���>g�2��Ln��i��������HνXݨ����j��F������S
���L��\ڎ^���8��JC5����]C��]r��<�Ι�����I��0aNVU �6������>��.�k��mŰ��ŵ���:)�e=���g0�4N�h\\�p4(a�������6tD"l$�k���<pC������4�Hz/�F@r��t������c/I����-;~�/�	y���b�ʩ#�8e�n�_r]SD	�p\84f��o�,�&��.&{M���r7?B��̑E�����x4E��I����r	L_Q���dh����
����O���b�~�_�/���'i���������wm۲�gZ�veYZ�����%�פx>����zX��LX�p1�<�n�𤃝��0�+f$]`T57A��Q�㥲��׷��'��1�vv��7���ȣ���2Aźۣ���W ��b�B 	cag��N%�:%�
H��M�bЇ�8�D~��8.�2(�Գ�5m���n��k+krc��һ���I
���h��;��DOr�m���+I'�n4�l:\,��t�7n��,��9�<'��������Ct�Qբ/�����AL �Mk=����t������3�V�oAjm�t�;Mynա�!�|<1fS�{Q��9Z�vq���:?�E�W`��qю�
)�;�-���ˇ>��r��Q�T�0�C�p���{��ǅ��`U�'��~T_*�%�����Cr�W�9�jۃ�BW�T���Oۜ�/,�I�/����5\N�aMy��.��TK�b=:(��c��>N����4#s�'�=�TM�CA� 7 1Ё�`C^���[��G�n"2Z��0�@9Ǆ�Z���l�Q�I�$�|@�H��i�؀m�9^�L���Q$#��Z�J΋����h߯�;59孉,��ڀq�`��>5�E�͛'ш~�H�[
#m(˿�R�-���r���:��͜�E�g���Q(��\�=��y��ٷOE'�K+�ޜ�W��q����L���s9��էQ��>��y������2qy�N���#���q10���������FQ���E7~ u!�Q@��u{�0c�(��W`p�-�ǯ5Ƣ��c�ї�}��xE�	�`��E�	�q4�E�JŇ�? 7�|r�B}:&b��(��/.o�;Q����4mK��7 ����zPN�!./��sy��W7۬�	�c�8����;�Gw�Nf����Ѝ�[�w>#�[��i$_�F��2�).h�5O\c(ZF}���Z�-+���C