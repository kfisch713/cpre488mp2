XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u����l8"��$ � 4Ѳ�����_�Ls����	/`s|TpƠ<$�	u���HD-��\b������쇤?*�ϭ�b �<c���CU���<}��i��vӷ�BO˭
Ҙ��ђ�{�j���A���a�
v>��Bu]$��O4i���Rs�k����|�Z�Ck;����Ի�̚���4VkTW�W�`��Y��Sv�Զb��S���ƺ*2}�oh�r"�kE,l�pU�|OK K �fmLp��Y����k(�=!\����O���t�c���m/��*Ѧ���NR@T(���=��Κj2���P>�?rs��G�O#��c�.�
[ �ӵY�GI���gx:O44^���
ܷ�Tn|gr��O-{�����3'�%D�=��@�h�U�O�8o��'(���z�Y��y�5�[����B8�R���	�E1%,-[�HSfԕh�8�Y-��r���?\�n��R�R:ɑsW�p'�.��R��5�P�?�@����ՃC�Xk��C�
Pc�"��+�h��P�2�����ݛ(�Ӕ�78wa<`��3c�e+�l:9O��8Xo5�U�p�>&��,�L�n𒒹�� H�ٌk8�X:��y?n�]��O�$���쀣�e�vq�z>���d	Gvf�?b�qu����O��z�l��J6e��VM	��M����\�����%@��i��O>܎�ܥ�2�KP����r��T�_v�Z���me���5�O.Zf�\3l����ȑ�$��XlxVHYEB    76a7    17c0
�V��ݐ�y�aV�����,\��U�$��J���4:8�'o�����^�6��F2��L;6�m+�q�x�3ѝ�t��D9�3E�ĳjv�� E`����T��WUG !�g;�A`�=���U#N�z��!�8��׆�ʶ��ԸsT��M8{���S�>2����ȓ65!�������@1@��[n��L=���٠;
�� E�� � U��A�4��l�8L�c�ػqT��1Ubeժ�b�+����m�p��US�!��--��/��l�X��%ɼ��X�R����^�cH���fj��=VW����{X�P�vt#4�^��q�~�e�N�}+~�(������P����]�	�)(��C�V�|��m��j�����h;��R���� Y��!^W�Ռ����8?C��˒
�J����zcAqpLT� ���e �xEc�J`����߰8Dx��c�ɒ�;(�y��XK��Ů��J$��&B��nW���}�G�{u��V4z��W�fX�5's�0	��!��[�l�EM����j~��l������9C�4Ͻ5cA5M�̯����<0!������i�ط��L�X��^L^�C�KYLʊJ8z3Ac�`A|���%�>��5��%�*�\:�3l�g�Ԡxzhq����)��d�����@W���9 �����j%uS�����Z۷F�F�m@8#���Z�s�!�]�߰]#A�@8�8�R�k	j��$���"ZP�B_L����4�;���N=�d�s�ZJ�0\۪���k�x[�����H����8^�Rxo���s�^�v���7�k/lf�dD�w�Z0![�ꁓ�>2<�Oy�D�6�2J���)*G��-�azO��� �v�mͼ�T��F���hl����t�#���3
I��M��j�g	�¡�����4�GVT-nh��5�X��G�@<?b�r�C���-5;a���e��y7��?��|�4\�}R\���Z���?��U���I��\04xpg���aI��v��4��~���)!�d�i�ɳ y���ߒ�3�Ӹ�G���s:�M�//
S65�1�k3��b~����UܮͥMV�����y
����HG���+���j<u����Lx�ƠĮ"�e���쏓Ow��_p~'�]�W�,���t6��.��0.!���	eIƨ�֓�������x��1�A�4��x֜Ŕ���k��]�<�{?h`,��`��n���Ƒ�?��|"(1�V�@I{7��}���:�;|x���kA�t��+�	}��N9� �쒄$�"	��xT͔�0��{IO��A����ݩ�9��"`���9�R�N.f�!����g�{���s�յ��@���� ݝo�e�n�t`�&��;�B������ރnB���F�c!������� ��*�<gq�E��aC�U1X YV��~�"ƑU�#~�gOg��pe��i<���,�n�Lze�-���3S�/�>��,�B'�\u������`��;��OF�K������#:5-h��(n���lDmt4���0��]��)3���p6Ḛ��4�i�2���R�Q�9�t�=-�N�`��'c��M�8l����Jd'u���Y��'k�
F�3:�6l(��
��I��	Z���&���'�1x*Y�f$q�v�|K;��	Xw����$�8[�Z��&gq�W�)��*�k�y'�P�������|��������� �3����q�y�1�����$BCR��ϻ�]���k�X#p���_ZB����7��]9*yx�q��x2O}F�}�E��:,�H>�x'��KE��{mY���� ���`�O5{~/��m����'YC�!	Z>_Rӑ)�
�T�I��
I6�%8�|�����4G���B^������{�K�����I)Uj~[w�O��ѥ-��|ی9b̂��}Y�����30�NTg��v	7�V�E�ꢴ����\Mt1郒
;[��e��3�B��j���}��"��������ı9_�Tf�M�n:�Xf�۳*2 �����r0�[�T�. m�@�Ի��)�1�D=��t|�Rm�z���&��	m�~�Z=1��Evz�XG3�\~�X3�<���mw��%9�٭���b勽i�;�9Q��$��A�=W{���#��V��$r��p4UY�������P�7�I�r(���A�����b&-�^����\E%��X+��^%����Bڨ�S�tXn��2�Cl#
�h����f��C씷I��L�������ι���	�nT�wQ��}��!̅�(B������Y��*e��W}�);�c�i�f�����Ї���������֝�}�l��XF̯���E�A���,���7��$��b�m������Y�c��x�In%xZiC�uy(t1�!
P(����³�
u6� 崁B� M�n�e~Z���%P�G"�jzdو�O��v~k��'���@1�=B�(�4 ���&ݜ��6EO7J����8zJ��蠠�Բ�X���=�*�|��P	&��S�!3*ms7G���y�q�(Ju�'Kj���3��U*�栥T���?w-,b�D|�Ξ+���_K�l��D�",t#6�|�R����a�L����7h��{�����U"��j�ߪK�eTl�k�^8*MLA�||Y����T�F�Yk�z�c/O$�ťrd㷱���Ú����Ե����(���Z:*aP1�í��&�z�dξl_���a�p*ڧ'�B}<:���>鉯��Q���5џI=��֊��e��pZ�	U��3���ZI��u�/r�Le�{%�H�(cFpu��;��"	H=���d�5mR�Y��*A�
��˳�O\}�Iʀ&�'-�ԯ`�0��_?�ƫg�>!uP:�w�����	���s��O���W��c�ZaV�ܬXx��q��	pn�(�<'�Puf?��8M���l3�,��s��%�`8�n���(~���E����'�F���?�Uf�;�-�߃9'�h�ynsLdk�bql�Ո�}٣�w�����eL�p�����qXM(�I�gq&8�A�dn�.�s��&/�444���Z� �˨�6xEr�F�1צ����2N&<�����rY����pv8ћ��:a7��7�3�Hc��uC�;��n��i��M��~^�v��2�d}m�!@��IˎJGn��z�z �p��h^[�N��|u���v�<|	J{���)�>|�igP�iAI'�3��S�	f(8�2�9S��|����>���Y}�]�y�Cc���0��q��~�'�hd�4�Fn�II�`���7��VIy�v���!>�m2��sA�"%�����ܡ���C�&q~U���U����y/�HX��7 o��"��9L�UK�	Ya!ƕ�7�?�G��7��q��,44i�A���!�3x��c㳚�ƈ5��Sr9����$T�?�66���������`-@rk�ԡ��}heCw��w��W���.�;�>���)<���^�7M��ɴ��:.0�l��x��zW�S�GZiUl��{�?9ia�rSh,f5Ir���k��O?z�6�tBn����y|Y�� �:�@6gH�Xpຉc�9�MxWNz_Q�J�r*��#�U���/�D��	v�v8�����M|����r��T�[K~�:M7��	�~u)����]����G;z��=J:��i ݞ�Z���f�Lj�x��`y���P��W"���^����8���5��n�߱�e/�ث����M�W����+��5<�W�Gy0�V���1����giS5�-�4f	�����f�g(v:�(�kg�ʫ�y5���i���t!��������h���}c�]N�IJ�6uZ^x=�o�:�� 9|+A9�3�y������q߄�̶����x��V���[u�[��6�����+`ħ�����Zx]��̲���c�u(=��H��F�́[#�9�x��:�q��fs�v%,�?0&jƉU�� 8����:��ES�n����������,�PN�2Դ����M����.����5]
���P�x�����P��.�klyw�E>��m�Z�� ��r�l��D�<���'����R���h��g��O��R\�����.�dН��wg����5Շ��g
�`e�/��:�eƆ��=9kn19!Lb�s�*���������a��r��p��2O��ףT;����2��6�� J��/s�y�aѓj�v�����4����ɀ)K��z�61S#���.��"�D[��CJ����ǁ�v��ӂ�C���<;%����Z؍qkU�,��YCN�*N��n�u��'>[�J�A�`���Sѩ�I�{a�։�� ��i�@�[��������EI�w���Z�d��fRӭ��L�����.�$P;�W�	��>?�=5_zMڞ���6d�ǣ+B}��e����������W��"cqS}.}n?����_}�e���r�k6[��N�i� �.���,�(y0w�i���P�l|�a=}�2�,i�ox���_:���Q��rg���l3�<��a�NJ���Tʣ��i.�E�M�E�z �AI�9uW�������J�T:�c����i�׎��<!�>2�	��������a�ܚ?3HR�b�M$�f(h@n�a�#��p�֧��rN�B I������~q�N��d���p{�;H�fT�Kk�O=���˒��_�䆷���9�O������C�/9_�E�MiX��B��x�^������\G�+��6��$�'�k�F]$.�׳�fX'��Y{�伄.Ὀ�P
 }6*y��".�ơ#�13��
2����W�E�̴���M¶�e���P0\٭��Cl?�3�C�K�I(ւK�ɲq���qޮ>�kW��ĩ�[B�7�.	N O� �^U(�xd秷�&�	ھ�|����*qN�}��B��`C0#j���ȗ~K�=o�ZFW�`]�_��&��S��a�z���Q>�O��<;P&��p��i]�9s�1Ѓ3�
';���\73�;�f��"���s�G���P]�y'���E����|������Ѕ���?n̆��`�4^6�q'=iJ5��u�W�8��oz�'~_�J�x��K�)}@�~���N���D�1=ZT�u��x���f{�'Z��?�~������1s�f1��f��,
���u���OS���B<O:$�������e�B�<��eu
 �SMIO�ref}��S3��C{�k�����Ҕ�3��;}h'��s�����.��Z��l��dn�w ݏ������$�(�Sba+6�7oG_L&IY�ɲ����G����:��o��טQ�1�)�RxE���0���Gbc�kBW�����TX����(�4
�!$r�F�׶�]b�_�n���9L�{��� Y�jV�n�����G��g%c�YPo�O��=BW�F�@��Z%X	k�(\4h-h��M`� M�-�X."ɂ�h�.�X1>i��O-�@f*�2{�æM._�Ni���0��mu�[�8��P�>\┫L#�\ƈi���b��0�2i�i�翊N�eN�R��찷����*4<�	�8�6}�1=��D���v� H�l����R@C�����<]�P_�#:��8��l���x�_�!�|��_@��1<�j�s;��M���<��5vx���Ф�#�j -s�8�h���s&Ia�������yhia#����_g��޵2G��"#�w�7����2���C�2�f���-O��8!����x6cU������Q߹�����(>�O��`�5�m���xǹpa�}�<���(\�E���{�rr���!}����K��@�����<P��I��Z&nA����X����������Y�w.�t,�G=Q�%x���37
���МJ�ɣ�