XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l1�*y9�FⅮ��3el�;z��2r��
Z�^�m_�w�*A�q'e��z���νE}�r���w�s�W/�nEp�_����˼5���3?�!��"�A��9�d�#��*i��D�����%�5%��<1)�
0j��T	g�V�����y�.8�B�(�|�#�B*<�/�'�v��/�Y���0u+XJ��2\7��@��A�@��V�S����털V��/b��t;1�jT�J��{ 
<���;�L��$!]�^��T��ZD�&E�r�5��߮,泄���c�P�/��,��Fg;��L�z�#�a+�JQ�#�u�qJ��S�A���
e.k� Ws�!Z��z�c��BjP櫾t�]�	�ط3̶�����߀��">p?'�����w���;
w�/���u������#Ԏ)L�p������w'׎���J�o��ǂ�1���'��|T��N��$����h��
׮\��ڞ0����]�m&#�|���:�}I����r5�u�bW^�E�hl�����u��\ ��sap��,Ў���@��U��?X�(K	��4���;�e�a����8O��3�E%�?���c?6'�Ǿ/��m~4ް��vާ#�'��u9qr�v�3AG���ׯ�{I���Rq�h������  �Ҏe!ƃo<����,س_5�4�,H��	ԏ����`tȆD+�?��k+!�e����t����4l/��.Υ���m��z�6�XlxVHYEB    5fea    1830��z�IV���8=�{��|�;�a��/�y(�4~��N�7��W
�a��T�ԅ�99,��a����m��}���F��[�֫>E�8T��-⊕1M���UH����>-M�J�#�_y2𦸣��L�e�f}��]�a�oegx���!q)��h��qW��C�i:H���D�P<�)N�H0�QV�N��G�@�5>�o��"�.�������Qq8�;�֚J�eN��	��u*�Ŵ��Z�� �[�����ϛ�es���b�(/jxnvoGHeɎs���1�Z�x�d�t�=Z�j�˲6�\z3��eo
��S�a	��}����S�BU�x����%kB�?��=��僌_����%�3�+����(Yh����%�b�A	Y�횸��y4yHW��p�#��Ek�Ѐh7g�5��^��	2���d�d5��1b:ߝ0Y�j�%a�z��$��_}�cF��>X&�J�������v�Xa.'����ɨr��oKBR�$���Ĺ��*j?��q
�&2/cF�E�}�)��\��׷����I�㍈B�_p��m�ZS�k+Hr,8J�һ�����9�_����
U���S�m��`���^L�v�C�p:��.v׷Bʂ�q�D��|Ve���MI����/ZW���P���@s`D|����Y�w@E!B,bi�j�r������՚6~��y�]e,Lf��1�)J��I����̬��	TƉ���'JUb4,�E�frf7��5߫���{�H[�}�E��?���G�v!�d����х�]{� �9��W[�lxsi"x�?���(G{�O�P;�H��Pe���KvGr��|�?M������)�B^��=�α�s�%z��}��d~���d�X��vn��wJ������(���=�G��)�D�r�w7D�������Z0tI�i5*ۉp�_�=a�qa���ޣ��/|Y��lgq罵�0TY|\�~�m�S-�Əo'S�:��x�H��=�"T�ꏾ.���އ�2|�B�$��{����K,�%� DR�4����ژz��3�ɳ�L�A�݉^���!�G��Zߥ�5�����}^^� �p)ʕwJE�j6ܮ�7o=�׋������٬�=&a���򖥃N��I��;(���֑W��8�s<0�*�P{'��k���O���Go� �fk�����(b��Ѥ��7��L3m(���*�:BCR~��Ì�_}�����/E�A����0&4���I�B���}���ߢぶ�-�D�)�=���&�����P<���'T�Z���ǨE���^!��@k��Vq�[����D����ƫ�g3k�!�ԡ�t:P��Q�M�1�<`��j�w�0����}�?#�$L��4���c8�d>Y"�0������eJ-4���Q�e!��Ɂ@r8�eB2��#�����tҋį�%��ڼ���8Ί@�o���\O�������f�"��`+��'i��Y��o��4Y��{"yknNL������)'T��㽩J�5�Ӿ+�e_�G�m�0�;]n�0Q�;�)�t�7��C���юμ�� rB��ˀ�>�2�/LJ��-^ᛵ�C�KQU������W.�k�]!��_��(z��JQÀ	��g*)�{鄽%�!�7�	�~���G��F�(��n�x�x\J�����1,
��E�����C��Ay�?Ib�f�c�!|�І�&���\O%�T����PX�!.�����~�ғ���w1g0X�ӽ��J����2�O�w��`� (���]�J����	�2�F7D�h���ȤyJd2Q_�������yN] �७��@���e�h1I<Ljf��� ��6���G���nT����ؔ��g���xh+�J����]��ڕYʸ�A�lx�⊣��1�S�9�/R�����3���A���D�raJq�\G���0��4�r6����|:e�!<�������P�E����Qo����~腷�KÐPIB�į�!��Z����j�+�n���ӣX���|�UW]���=�ㄯo�J���s�N������ӽ����j/|��k��+0��y��"���$|+�T�!]�,���*}�k���Җ�0bC�[ܯ��Mdm2�]�[�'��k}�ʑ!�����Њ��'���y�xBK�C�#l��\�5"���oՍ�JHoz�t�[�ą������{�Q�P�ڦ3�up��$���F~o:�N/�Ia,��Rÿ?��� ��)��_�+��S�	�/N��]}�����Oڰo�C%���� o���:��a�	N੹�S��U;���_FET4۝[_��Wk)���\C�rx��[)|1�,�N���oo�����-|PjK.Ql���r��(b��+��n|��PV��z�>á�r#"�r�9��ɰT�/�B�"	߳����JE�Qe��vԛ��{���=$[WKT�	�2�Ӕ��Cqne�3[&:[�7S�"61���/��&#l�����au�?�#r�B&���L�|�9N��^��[C2E�TyvN~�;�Ź-�76+��}�xo15�t�{*�6ր��u�(.bg�v���
P��p���+�I4�w���kc��Ǎ�M�L�;�ê�g!O��i��wE��ٵv5o�ӛ��q�J���[[i�$�%�=53.:6�z���!�܆�6Ɲ�Ao"��Q#3��ۃ�Z�����`m�_`g&�-��|M� ��⿍B�aB�nz{!4�s!*�yB4�X��t��%��[��"ɲ �,Q�	����!�F�D�# �4���C�m���y0Lb���	�Ĕ�0n�)���U������:����D�d�1#��H��vw3�2�V	̓²�퍬���r�K	pM������sq��Eu�;#�����l;KM��廛���� >R�T'��<i�緆2�d���������=A�ZiI�����?V��%��j������Fy�&f����f��̔��6�?�kdjP�m�#�~�҂Y�f��!g�[-.��F�d�r$�)^����Ze�}&r����dǄ#�
�w1&�I��[�
5j����gQ��'�,�~���G�0��1z>#�l��j���I�����nz��"��b��RH[e�!�,�FOE����xt
���/3rp�	c�D�q��щ�]�3���7SzV����I�s*㕗�B�:�����̿8����-� �['����O�AƢ^��S��֒D���e9fu�W���ӳ���!������B+��`Ն�*�sq�G�"��y���v<��`秳�3� ���(F�A�\���L�;7mx���m�����K�����p��V�LYO�5W3w��q%Y��=��$���B6Yo�X�@Ս�Q;+	�vJ�M�c
`�V>�(�+G+/(�*^�Z�P�t��D⛬X_)dx�:v� �QM�o��x�;ئ`nxj�����̿��/W��(���BC�BYxaB�e_r8��E���.����@\[�r]����"������؍FG��aMx��5fM����{�<��ÐF�O��ds�ܶ����^ǡI}t�.��j�cI�I��J�;����֗��0c�����ohQF�:���4}��[���O��0�#�%Ǳ>�wy�zxH�������bg�������{�H�{������Z���X��ā`����͝� TW-[k������N].Ŋ2�4������{)+��1��AKp����������Ο����qK��U��(���xNN�<A�O���b;�|�h��J'&O!ʤ�h߆v�>һε-�?���ؕ��~|�*��;$�1�|k3[ZTM-�_��"�p��.��7W6�|B	
,�dd���^����+��E�\�����A0h�#�i����C,u�˓�K`&wd��$܀7SQ�55��:x���[���"ݍ
A�4�W쳦F��}�pd��6dJY�/�]�X��?5��j��P���Մ��ޓ=xKoy`�G-�>3�25w�eD��9';ٵc����Aʾ�)�Q�`���h��	��L�t�=�#1� ם���y�\_��/�����ӡR�lY.=��?�{jХ��-t=�R�w��B�0�X@�3
?�����a�+����fw�.!+���]������X� vҟ��0�?�{n/��̳�.]y�4���Æ��v���F�����,a�R<]̯��2x�pJb7q�K4S�7wya�����$b�w���I��h`��/*�N��o�M�.s����uo>m���	����(�������Eh�M�]7�����V�o�ـ�E�����v���(���#t���ɎH�fy4Y�[K�,���z]�
7@vsð���C�� �]���L��>��s$�������� �|�ׁ(#�׬zu������̝�(�k�G�@L(��n@8����㓚ķ<〖>:lc��ȇ�o�TK�l[� ��*4`�-ma�W8�6Ԭ臐����(ޜ�:��s��ր��d}Ýk0N�V��"(�}�U��M��%7�� �N�q����C�G�����Z�u�xcc�~��'������2Sg:ekX_�u�(��ʑ��ہ2X�^_��d.ʐ?R��w�f��y��jQ��V��^�\��4G�7�L��h�[#X�1F�¸�]�S��5�����'�M�VB��Åi[�1�Ʌ��!��,簿U�Cbٿ	��:�O�ٽdh��{��ڄ����s�h��m�{��q
���!�[\)pn,�F�{y���\g��D�a�5��*Ϙ^�����b�=��Q@\�Fc��nj���y��it��?Vd�I���C{EK�t���t��C�¯��G�7尷���n�-5v��2k�`��Ѱ��vʂJ�ٌS�.	2���yp�=�zqp`b�H3�Ɨ�<u�K�H�My�ԞD���K���Ӳ�tQń��R��S G��ի�D[R;C���.��
g�Н�w_<�R�=��@^4�D�ZH`��T�c(�)��,{�~ہg�h1�IE5�n�G:�|��䤶qu*�]���{��O���xy�JѤW���J�V��Z����ʨv����%���V�&I�x�^��|��8"o���fMfxg/���h�vY*`���R��W�:�kd�c���N-�[�P�x�FJ�*["=�p��$��sh�/�)��=�.x*�S�9V�a���R����ֆF4�5���E����M��F�C��m���Զ��7��������_|��|�d��C����*/{��x���l<Q� ���MЮpa��5"��gם�>d��N��|(V�OmƓ�����
���Q�#�'6aíB'�T�
|=��\��<Y��o-Ջ�^��xy3:�,}Wa�\`	���Q��o@��s���p%��{��vw5Φm��:Ȕ-�b�_L�6l,��L>K,pj�(���
��d���l��3\C�d�e������v���-�HNw�7��Ły�����&\�V�Q#b���h�U��3m�w2(��n"|,�oa��&I�2+��`������b}�^�B8 �I&<;IU@U�++���տ}[5��	~�Ι�w�֚;R|R	L������\2����.y\��>�S�G��ΚOaP��~��U��)��c���N�l��SlU;W��'~�30�(�'�UD4R}�e��Mj�o���hNeL�I� ���}�t��6��k2���9��{�9���({
)�'âun��B��sf�E�c�l���9�v��
��e�z��LD[��~;hS��d|�}�l_xp����ˡ=�SM�������	�)H��=Y�UqVj��R:��TL�Mh�:�7�����׺�z=�=J������[��i�"���$R���e�6�ٜ�%�9�3�-x}Jઇ�q�r lwG�+�v���6y���fY{>�n���G�W��

��x���f2`�<n9M;i[5�T�
��~��+7�/R
浳��X���1�ub�f{b߲/2ɨ���tQK��d�������`oj��̓]��Һ�rc�&5�����Gc ��[K