XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_�ř�KO�xޙ���R%�ƤzjW~���G�p.��DV�@�p���^�Z@t%ˊ��D&�[�'�����}^�]9L���70�ńZC���l���=瘨�J��O_~��U5���Z��*��o6���XY�c�5�@v�q�=�E��a}Ƿ�\c	MG�:/ !�`�lY��>��7іN�����[TyE��S��:����)�퇟�$�<2g M��&_��%H�e9 ��Zb���}4l�=�� ��7[ꍮ�1
P��r7���
��+]��{(mZ�!�価ڛ�˲JD�AO�L��Y3�ekv漈���yx� ����RÛ�p}s�UUWG�f�� ��*&���y����l�-X�}�^�^<%�YZJ��w�H��岷����o��v+P�=��]L��6GT� kIi&���s�1W�C��W���D)�n\�"%�u#�q�R�k
K�GIf:��p4��N�B�dsVv��4�i�J^���L�p��TIL>`:��쾄��'��Ǽ��9�y��e���u�,�G�<J���A�9EM|�Y����`�noDJ���<�b������=c��_���J�Ƅ����=PJoE�ʛ�MT"�Ü�Sۯ$q%��+pGԫe�:7�&7�����!1ňU����	qr6g���t9��"��>�S"��_�¶T{ɡʄ�`X@U�[.��ƶ�!+b���yխ�m�R Ēd�Z��5��_l��h�C�asPŇ����XlxVHYEB    da59    2e30���'�$B3�<���W�أ���.̦8�O���ĮԈ�L\��?�=}_�������*{�h>:�dA��W}��.���#�iwL�.�~�����4�QG��k]W,�1�!���hcC�h^�����'�>7��D���dr�������d_��l���$\
S.N�-C8��Q�Cd�W�fy��5@�ꅔ��\B� � l�}�(o)q�y�'�V�[d#S��$$w��D�0�I��k��uݠ�X1kf[@��O�{������*ʕHkB�3����K�g� �ޏ�e:�|���4�1_��`B�#�����LV�{����OHְ�{"D�V��k	
�i�n7��Ʊ�+R�N�{>��=����`�"�h�)����O=��H�-4F~�y�(l����9��2vә$�Q�fR;��NT7����^T6b;�&�E$p����P��������oa�Ƒ01n[!9�;��Z҈�3�H5��Q�����w�U��l|%�,�Ek=(3��F��U?���6e�Fc-F��@p��W�m��+��V��٪x���Y��thFE��+�p��pN��&�S�Zq��>eO�O.&��� ��0���M��H�u"��?�H�-��0�2bꑙ��IǄ����OR�<'4�3�8�5��E�@6̆+��PH���uK>|I7FG]����4�jX��YaNbe�z^c���OL�
��I]�Jb�f�6�g��cI]'�;x�o{V�Kْ..��ԑ��0.Nc��_��h�#�Ԅ��g�nz3�j��R��%ͥ��e�D:`BS�
04����g��w"��ûL�5
���`EA���ud��r\��W"劗p��G)��%����*�Q(�eYKi��Z�n��j����uB 'd����H9�WLIﻛ����4)�[�^Z�u|���h�҃RǷ?�0� VD�Q4�utQ?���o@�=��]�q���V��	n{���
�:��s��r<ܦR���ʪ��}=��H S�*.��o>� +'�J�xX};"��m�R_n���j*��ސ��ؼrA�"�Y.�%�n���D�I�<��2��n��mN?��׽f��FL[�E�z�-�&�C��XQ�/�������M�.-���f�M�7-�%�׹/pQ�nv�6�$\0�O��o�ì��\`�A�U�r�(%sS���m�N���]Ծ�%�GpUV���L�������|w:����z�e�]��zA���q��d�����}��T��4[�	��|�Y)�ntY�c�(���~��yyΎ��`]!W�P�"�4�v��ք��_���G� ϋ�*7m�W���s�=��i^��p��C�ZS~�ܟ���4�^��Ӧ�Tf�g}A"�ŷ9؛T�#���;��F�.8;�S_�P��'W�}=D� ؍#�׈��.Ь��-&���&�<��<*1�)�$jQ"LK�s��7TT�Qw!� zC;d��ޏXBs�1�f��~w���a;�'\*�MY�Jj�@�3�%�d��}�#U'�ɢ6| T����D�٦^��Ӈ�IΠ��U�!�[���n���p�]��U
?�ו��JH�W�"Cy��W��K��u�������▹/f�k��jibX���6@��i��%�����v�m�?�1�y�392U��n���S=f}��n3����4��H4�
ʃ��I�E�JϮ��uD���VH_9z%i��	�-�/��9
����7B��n����siY	��nG�xUO��OV��6k�W"5أbr���� ��9JЎ���Z�=Z�8��li �=}��I�A뭸C`�o"Z���x�a�-ҼX�hm̂�V'H�xo�ץ�8��N��,PL��b5t#���?X��&��x]:Hg)�����ᄯ��9���e��\"7�]}'�;��	WM��E�xgZ������N=Wup�'O�5�3�i$~�V�ݻ�mU`V�(�e���j�t��~�U�'����1�%�cf��rl��z�c��A|��UK�v�".C�'K�j��ӟ��Ņ��K\�q�}'3�!�2���l�ꟍ��]����)�&�ς%�E���� X�� I���?wej��w_i���ū����7��9��	�s���,k�:�� ��D�U��V��m���i��RU��S��]l��T���C8�E���M�Y�����X��F��m����Wp�z�T���֊25���[F<���k�W��~^!�Untw�P�S2J��Q[��x���d"��l��9|��LՀ3����2V���.j�O#����/'^�ܣo#xd5ݪɭ�j��ȭC��Ř�W��C,m�!;�9���{�F�#nY��z�������Ⴣz9,X>�]x)��m�*��?'~��Ȟ�@[�8@�A��|��O�mD��	�T��\�Pٛk���j���r�����+��WM���;����%��H��*��=��tul߹b(@0^l���S3���J^GR �z�+����[4ޫLjU�&��U��3/L�3[�wG�&!o�;�j6�tȲ"�]R ��@���L�J	!�0[�a?���(�H���+2�K��c�z
�TG�=��
|���| [!w���<��^j#,pTܐ��l[A�[�Ɇ�����&!^ M���9A*�j�\�շ�:��||�=j?_}j��#3�}���+59��ô���+Bp��=5��S0�]H�a��$��y�땅��q�<u����X|��AG�
��Z�v�SHsbfI�#6|c�x��$ͪu;�CW���� �ꠑ-���vGk!t�r�O�9�i>��F�(�x��¶�o�8Z��߫��lX*.���U��bTt��EP�BeVpN}+q�1w�4�X�F������b�����M�� ؠF���O9�6��jk-� �R ��o�/8��bqA9��'nD�Av`�.�I�Ɏ�>j��o.h�M3�B�m��]��xK̜Q F,�%z�����?/�B�+қ���Z£���u��33�g���}9�L��W4W˨G�2�'�m�x�	ڎY�[�@�5�3�"ǫi)��=��N�ؖyKp�����}����~H��%��D�f�q��N�
���I��	eP]�ރ�F��b(-A�t ��#i%�J�M�ƴ 5k�qj�=���H)��L�9ʵ����'	�P>|}�u�սA�(���A�sL����]�[G�a�n9Ԯ3�&��=	�]��G�v�*֪~����Ly����a2���E�1oݢ:�60���E��Es���p���ӈQ�1lء����ozoj&��'P�J��(�p��^[@]��r�} ����:*����o��'
���jN�iZ�چlM��w�=+�Xuβ���bg��d&�pP��Z��J٤6�t�Шm�!��7�!���Z���2�@~�$��2[G7^v���U�6���m�ER�M�T�z�Sn��)���3�"H���;E�nj�cT
_�]˵���֢�m��#P��VA�1g�����8&�~��C��*����C� �j�CB��d�J�
j���o15/�ڤ��|�S1�aB�U�9�bŶB�Ӎx���fWϭ)̅{��]�i%)k`�M��7.^�.��{�-�4c����������aOV�2�d��=^WA�M�{��������H��]6]���C.���מ�ŽK�-���oS�i��e{�T�X3����4h�K���v�G+�j���oj/�~����~��c@�<����W�O:Io6$ Y8�|����'A����֗7�^F��S��8�sͳ�q���T��_�mz�_�0�h^6m����o�b��.��T��x;�%��;��=	���h����SG��@Ԟ"����Fai�6�Dّ1[�Q�mZ���Vu�`�E����W�u���a�N�{W��+����o;�M٘F�,�˙(� �H�/�|��`b�"C߸�F�2�Pb7<1z�
w�N���B�:0O)$*)��L�x����~�t���[kV6�*��߻�s����� J�˵Z
�����L���Yo�פt�w��+�yг��-�v�'d]����΀�P��rZϚ+y��:�V�ɼxj����I�(r���<K�&�Q&)UY.c�F�v_܈�C����T�G��ص�<FW"�;��T�}����Mt03�/�L���S_���`k�및vl<�� �*>�x���a�k��^k?� �n�p9��gܛ������S�:�e�Fe��E.��X�7�>ߍc�b�4��?�֒g��܍�㶶#�>A�?�v�������������辮�]�@�<h��`��t������1z��������Y*����r��ېɊ-u� U���g��h%��d[_��Y����+vt�H�e������ӈ�[�ܩ���[�q]������~R�<L�C���_���qc���R/M�*��{�Z��O�?+B�<BE[����1�_�.�]J�k0�]�oH��c�2�z�I�Ł��$!��7��^tc��O�f��n!�n�,U�����CEp��oRIʖ�Z���c�
�����cB.��%��uJ�ѳF+�4WhǺ�Z�\/T��}�a΃�c)҆�$��=z��`�IC��}��Mr��?)�l>�~nˍ��JK��$��s����f��d�'k��`�)�J`��_=V��/�f����R�<�	͚S�㤛w����up��k��~�F�z:IBf�Qm5��"8��Jv����t��^bΈٞ4�����Ѐ�O��b1���\��k���1Cg�|��-�����ʈs<B� &%7A���R�mx5��9�������b��'ڔi�pz�r����N_͹厱�*>/=�u���Y��G^��O�W��I�p�A�Y<5�Ѓє� ��Q���&��ϵ@��ha�ߙm�.Y��i�8�0��i�O�+��ݑ�4��g�W@���;�n���#cM� �)q!9�ޅT�A�I-6��| ��]�ͽ) ��MEK�|]��t��Fr$�u�,E�y�f�Pb��[��M��y�Ele�~�X���B38]ƛ�����~�B�	��&d��{"̤�Y�.�eJ�kM�I~C&��Bf����PK��Ό(���t�}^�֌���Z����c��;́#����@�SBwOZ�Q]$������<��
kS.6;�X[2�r3^��Q?�5��o@� ~�N��6�9�k$Z�o]�l�� ��SD�6;���\�Sgi�M.�E'�Kc2���a�M��0��W87��AP<D��1�x��]q�X ��K1L�!�2����J���ky��+�Q�����u�﫮�G���e2+爋�u��B:8P�;3�����`���w�ๆ��R/Ͳr�$��J(>T���7f����B���o'� ���+7r^�y%�v�B�A<)C7p�fi�m<y�����|9���E�1<vS{�;��]�x��\���7J�eV�k[L(��
FF%saF�ꥢZ�ڭP��%��D���k&>U\�4�  ���:�"�h�EJ���T�.@�LEy5��1���B�A�~��K���t�}H,f]��5�Al)���d ��2��9��FծV� ڂ���h��Q����f�	D�0�&A��1�ŵ��un����o���UW�"�����h�mk�؛%��uN;�O�ɇ�.�!��*�iQ�,��A������^~u^D6��,����z���xx�y�q���f�'ɖb6"����<χkJ5�]彝�֧V	���.����+�ϙ�>�.�L\#��l��׋��'C�����(Z���4��I�j�hƆ��0���p�G���U<��D����P�����*��e?�D�d�[����\�En�}n��n�o��$����;�?�V⌣4��)(yj�ďxz�R�S�vjIC++𨋥%^���'�N�L��;>�
�SE�jZ��@�^����u��
?�L�S}$K�ˤ\�j##�}�I�o���Y�
����	�8������^:"�=��q��p(H�Y�;�6�����,(q��'F�j`�<��c����rB\��ɢ[ D�Rk��A��"�a��Q"��'!��XHo�12��sTYc7fL���cki�Ջ�{;Ά=>xs�p���I�|��j���:��=|�0uty�<�e��JE'AJ[vt��������ueb�XP~St˸��ѷ%F�AM� ����d�7lpt�|�v�v;���6E�|�PZ�d�]�^C�7�u���$0v�U'��÷FW_E3�.�M�څ/�=�&Ķz���y��څj�~V~l.1 �|g�����5ZM�����qD��`�q�8i��r����EK���w�{b2�JFY<�n"J�hG8�d#�f���~�2��f�+��*p#��76�LY��FƧH����|H�:~�t�F	F�稍�M
�K]���YuC#zzLgq�r�<aZy�
Sʞɑ㠈�LL:F1�İ��U�:��s���e�K����/3̿��MnY�eY�]�@q��-u�~��&]!t����u����J|\�����u�(Zb{���٣�i��>Ǉ��1`��z	���ţ���G��E֠q�> p�F���[�--�l�/���+����9^���F�
�s\`��[�<+�=�0˄���%�{;
�O�[1x�7e��c��I��(=,`�9ٌ���[}{
��"�w[�1a���6�χ�DS��A�<@��&� �cxTO;H`������|�Z�97�S�����r"d=��߭�G����E2~�Y��L��؜;B>�sH�D�c�5+'��U����Hw���X�������BG�k����l�d2P�N�I�Y��������E��
2�����Z�W�H۶¶���\}:�6����l���5��f�E�G��֭h��-�� N&�D�r*�D�V�m7�p���~khw�^��M�-t�	��	`��y�D�{R�όq�2�F#�&�^c���G����oWi??��L Q)a)���[>�`?�����w���؁�f��Z�W�ﱘ�_ũ���ؙzKt�!�\��oʧ��yH�Z"���g�L`���(M�o�4p�]�࣑x8{Vgk�c�� �L<?�n��7�~Zf8GEq����?fc``*;@�5'�oBרq�@(�m�mPs��M;��?s�{������]=���*�R!�D��0N��B�$����?�z{0�Od�'���Ǵ�v����	m� 
���v�O���w?��&:*@���F�mi]�c" ���fh�m~�>t嵂����(�����!�AXχ.���we���+�c��C<}o�}��v􈆾۞x��_��B*L!�����$lbk�`};���;��>X�2��1���WU���"��j۵8gx�B�*��_�xCD?t`=\�	�  ᯤst���۞r`�"��� (���s�9�l(��r��#����N� D�~kg�BFR��b�6K�+������D5(�f�`�б��pspaW�C���ه��w�������t�?�.
���,�<��X��׋C*	�7�pa��a��Mc�������ІMve92��͍`��b� E�D@��U�3�x��uB�ͱ�����j�L>֫Jxԝ�$E�a�ܭތ3u�[���݌w��,]QW%e+��2~S=�3~ր���xz�miD��O�E�@�2����v���ۅ_��V%�7�zҷ;	l��>�p35ݙ�i���e��	y*�	����Xx11�ȘBㆽ���0�̔mP���@�?{���g�����r����˷-�XI�=A�S:/H��C�`%�#�� j����qg�mvC�7�۬�����ů�����B9��Z��]�eĘ�ގV��uA$���y�o .�[���� p���[ȵ�o���ヮ�| �l�"�3�|.�&(GJ�9k�2\�؆���21�B"�D�i�>IG��h���֏��I����U[bu\����jN)��	]��(Mm@�[�=cװ�Y���ʧ���t�m�fwjG�+�k�lK�b����c[Iӵ/��ʜ����B��+���vM7j*�|��x[���Tf��g�0��7fm8�0�i�����Y�ƈ���nS��.�SRg�*��̙G9W�[uMC�4 ߟ�� ��&�Q�̀	 *���7�<#��3Z4I7%�I�����$`Z�_U����f�����O�i�Nu?���H��fb�cPn�ZgZ&=L�Ú"��(�g!,j��z��`Q����
�R��=-W�T�v�za��	����]�D3�w�8�+(J�F�O�2)wB�� !aC2����m��؈��Ϻ秠D�8���>g9��&Tc�8�N0���2�n�5�4|��]/���l��M� $nB�C=�o�  X���[dl�M&�JZ�D�
�":�N~��{��= yI�)71�W�f�U���P�c7��aSc.�֎{�%��P��O:ݬB����F�qs���JJ~�@ǁI���T��������Y�ud��T�"i����~��A���6��A�R�T\��'d[YHL=�|��5�^���${��b,�?���ft��娷��UlL<��c���nՀ}`�A�x@��,�!Y�"���Hv�~b口耥|.�o]򏹉kH�V(,/�q �7;Ÿ\_�:��k����s	b�1e}($����®����c|�`�wp=B �.;}{e�%�d����y�CdB5li��JR��|��3�6�%?�g[c=�A]س=�~������zR��N�+xp�Zڪ&G��ԥZ^��5�}�Gf�8d��>�"?��+T���B�=�V#J���g	(�u���QF.�O��;�r������\w�Ja�?n�Y x�u,�4�{���YV�9j�e_��1�7�[!�Lq=��a�|Q��� ^�{IpQa$o�\Xǖ�����x�����m n�\8��BI��W�K�T�?Y���(���)�%u����~�{غ�����jցƀ�6h�[P,����Z��	_�3�o�mv�āz�w�<`�Gu��pF#1s�k4�|
:t& x��-X��JW2,M��r�pHG�I*  ,�39Y�ѯ,��9.�ڢI��)*�N�u��b���՗䳍l��q%��Y�?q$v^�~���O�1��$��;lo̹h�i4��{�eP�'n˘�»ӗ� m�nS��?�N���C�z�:�JD�7����*@� b��W�^,���s���PӸ�4�A�>�7(��^K]˝K�����/�q"ZM���9��i��G++��#,odO�n������Ӧ�%�)&�ԟÂ����qN���
s�lǅ���S.m��{X�U��͸�H�q%!�c���V7;\�N<�dX.$��R��������6<��peb�b48�����Ҏ�EѧQ�m�7a|�jƘ��%�������+���=,:䔒j�]�P��>��W��(�.p}cc&��	��Y�j�12}��E��a�7��f�#�C!�|��[���#���4_O���~~	��G�x��b_z����D���o��m�Z�yas%�v�,��_#+d��i�j�oz"��L�8���7�N��f�&|��!A�f@ ��8�v���[�����4��i��
����I:=Y<���R�~_��cD�t�fQ��>��
�e�cV��BG�K"���%�$��Qty�h8�نB�58
?gx?����}�g	��!�s^7N��5w���PWϧ�)�l�82��25�c����o6~1DY@U�X�b�`?8���}��������I���@m8{�j�q5����ﵩ�RΡ����Ǚ����4�
��`Ñ�[AbC\�h���b9wև�����=��%u�y�1���4���4G��d���5�. �ڸ�����+�,�ɵ��m����?�kEx������T0]�җNăW�҆���ش"� �e��Ӽ���ʿ&�v�P�,����l�0�A���ڂ���v�����1�^-r1�{v� �x�G�dօ�&��Ƞ9R/,,F�i���~ջ���7� ��>�	�P�<[m� x�ֽ	���!��ء�p��;t�-&x?��4�ʺ��*��L�+������	1I��o��Ҭ�"l| ,��)Q�ay��R�Y�!��.���������[^�fAc_��n�Z�rl�ϕ���}b\	3$#;%Gg?i?5�$�0/���2��D\5Eu.��o��e��E��h(��߹)�0!�J�f�wl='�6ѳU����:MD�D{�:�'QM){X������i>�y���>E��y�&q ?�%	 �$j��/d��p�"� ��n�Ow�l ���'�n�'��Y)t6�^O�Բ�`R*@X*o`L>~�|l�w]����F�q�G�]W���!�ⱞ�ow"i����o�D��?��ƶ˰�q�︲�I��g�1�ܯ���nt���[��(�:	O7���$�𹛊|�%Ou_!N����XD�����ġ촒�[�>�et9鍏��^Ֆ�9T}�����l��Lv��Y�b,:�����x=?��Ϋ�����&7`g�]������͆�F�A:H�?�0B��<�����xf�7�goj�Z�9����@Dν�<�����9xB��+ ���Y ��s=޸P@r1"�E��@�����}n�/��Kg�+.��F�|;/�֛�Y6��>;g6�ֵ?�e�X�$Z�<�q�T�x��6�;|�JS�� '����)�XxU�D1$�)��x	s��$���?���\$�߯t6�o��co.K~�,/�T�������/T��.��t�Gb)7�I4v��"a�������r��3�+悮����G�ۮ$҈�$�rE8����,¤������\�e�e�;�"ʇ��YԮLo�}ۅ�F�*�� ���=r�	s��f7~~7�̿�*\��j����>���%�G�;;f&�5�W��V��A	Y�%�������cA�w
�ūv�ǚ� ў���O�x?��Ց�:���O�MX�ԣ�I�4Ӈ�V�F�`����J)�:�{�����	Z��0~�5�C�F&�Ŕ�(��pb3[H��_t��*�eA�j2e���@�E�s�]�(�qgi��������Cw�0�D��9�mbwv�Ec�{���v�3]`�%�����m6��}�/��굹�T��7Sn*��G������?p�ᥱ��,<��耶�	!_���.�T]����1�T<�DH���{���|�a�"�C�RAA���<ǨrC{F�d�8�Gf��*yp�Gz�����(�;�)X����n6�sv�ҙ@qN>{��	����r���";4��%e������e�ݭ��Dk�0Yi쮌�P��PB9����[�aoГ;@�P3��v�)��T�E�@]���8�l��W�����7�`��R���ݭz�3��c���I|�Jw�/�L���N�󽣏�5��#�dC��-pv�[��:P0�R��3��M�SwչS�SFZ9�JbƓ;���WePf�*tYI��@x�ϰ�-��N���Ba�p`�<�'���yI��w~�)#�l�#�&�P/��=�ۥ�J�9�