XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n]o�s��d� $R=�Jɿ�Ⱥ��#�����2�Q[@����7��獡3��� }�rKX�WL�_���(EV��M�S���ɫ��z�ew�����3lT�`b�P�3@�I*r�_��c;ڞP=\���K�u�'zM��d}*2�P�a��$��1w�2��1@fg	��u����2����-�ߥ�"��G�ڲ�L�n#]�.;|�k�[aO��}C\k��ɴ����%6�r������=O��bm �o6Pk8�,����9��!q��������Y�q�'�s�à�E�O]{�,��⥡�C "zSB��mS�ġ�T�ǔ=,v��q����!8��Z4���Q0��(!����ߑ\�c��0�-j<x�S ��+X6�(`L��L����O�3��|类�у��V��b��W����Lz�"���kqS[���Y�I���U\w� ��NeI���������ȑ9�쾔ऱ���-�&%���=��P�o�U�Z�*A�w����3	��22��X��[[��xc��C����e]K�߁	�d��P���m����A��\Kr7�:(4g/��_��/���[q_�I��|��:)#Ʀ��#�š��A�lR��~���ĭ[�MW\��r���]�k�;����5BY�J'{�*gUp�8w$3AP����G��2����ͫ�����)i��-BٴW�?CTpy���1ya|i�T���r��6�b�W�W�2b����b���^{�@q��P��8� �6XlxVHYEB    17d8     890�RYȝ��L�t'LG����2hH�BEx� ��8��f��6���~3�������t��#E7H\�K�dj;�զx$Y����W�46�K�Y~2�S戵�H��}��SW�w|t���J�����@P�9��bҵ���XP9���e�J�Z �kz�1�qH<��S�I8����fq/c�	��c>ׂT�
��Kk����,�h�I�\��r�舔hr��THu���ƹ�7M���P��L;�O�Ӹ��Dt���l[�Y�Dji�p�����IX��At�Rm���|���)���Y�1�]�T��e�{Ơ��~/wU���5V	}��5ieC�.Ğ�e��O� [y>��J�5���Ͱ�0�a���0���������,`�߁V#Ti?^x�1���zlEk�~�w�+���ЪΊ�T2���;�y֐�Ƕ�>�p輕8��C �م����.�}�t����1�;�Iw�M*�DG��%�=<$�fDf��*�9�G�'��q[
�f��M�o������ģ��j3��!2Mjj=�:º��j�.� |�����u�zR鵥N��,K��}[5?@'�>K�ߙ"�>�{S"s���A��<O#��u��9(�`˿�n,�g�S�8.ϵ�  �>�o=ꭳ�}��8���~x.�����^�����2�SݚȌe��h���b]{}QM��?e����`Z�q:�Ek�
*�@��pb�F��W��>'�. ���7�\j,�
%|�,�9�olF��
��.`$r�E$QV�%&Kϫ$1�$^g�{|^4�h������(��$Ir��]�N��܉q�o���rh����'��h# ��r>3�}C��X+���)�%�2û��^ U��<�B)�� �)i�8��ׯ:����JMs�ޖ�_�gjk:w��gM���`	D;G6�>t�6����i�q�A��dqݨl��k@a��#��`�q��̈{2݄FM9 ́����f%�0*�^�pv�:w��um��=ɾ� F@k�jgY��G4e+pb�Gr����!Τ�E�Å� y��I�܇N_<�5��ܼ����pz��*�s�d�CnF���?ngL�N���<N���ks�gݴ�%?�W��(�Ը��֬^h� �\�=�\I���!c%`���U��S`�T�N6_G&@.ޙ��֜��H.<����uqa���P��+���;O�����K�7�NjU^xK`�X�X��D���_�\�.`|'./�,S@�0Fg�$+��<�==���{��O~,�\.�b�;��F�h���,��P���B*�9��4�y���b狥Y���h��$N�c%�%���QG9��R��{�m�V��$���]��|��z3�j�y����PR$i�S~ڦ]#3%R-+Y/�ow�X}��ڝI:�+�5��g7�H9UT٥)�!�C�A��$�EϽ��%�M�w-��o܀�қ��F����e����^��|YZg�N��&�ly�]ƍw"[Zv��Xô�o��iq��Qk>1@�eK"���P縑�/��<��1��ˍ.��.����SgF��Y�b`�>��{�_�׆k>�^<��< �@�~=�(���lL"#��N�����cO�v�|�7��r�J��Z��f��������
�f����֍K�ؘh�
��x뀢��Z��{��v.���M�"24�;��ү��i�A� �{0O�� 7J>�o-����Re�M2+�@���1vO�f�x�[�bl��Q�� ����;��#���%���<��_���
�������x�CsģĘ�f���_L�]�೨�Ɵ�J�M�����$�4Q����n���	K�T�Q�c�x5`��1Jq�?�}���Og�#������C�O��:�������00�V^s2WԂG�0�&Us����c��Z���-�I|��Iqԋ�����@J"l+��B����!�l"~��~�:�R��#?���h$��^&�l#���)+��F���a�6�^%Y����mﭽ���A	E�nZ��+��E]n��k	��x���@��f:�)m�S��QSV$8Ϊ�"�1�kg;��@�9s{���]�n��!�[�����j���*� +�C:�w��)ώ���(��B�����o�#��t�`f��