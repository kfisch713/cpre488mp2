XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��EF�X�o&E��(�z}�T�?fh�V�~�G~��G�(���p�@f�[TѩD�n���gA��v�Z��X�Ω걳c9W�Տw5�����Y@���i�k8}�}#���	���t{�2](W>X�/±_�%e���>Ǟ(G����1u�Xm>H�KkYX���"�i1� �3~1A��R�����T���;Y2j��vCg.4@Z���]Ցi���ғ�T����(>1e�k�ۍ���Sb6���רXZL3r���oԕ�vn�q���m2��8-@E��� �4��tm�s�A�s�jiv����}GF	���a�߷µ�)��9�����R��@t�b�3�;Bs��x��9�V"�Sf�L��slbd���.S���	��� ��� �e��P`�?3b[�۝��zhˈؘt�u'E�W�I#zOB	P0��l}�~\���a珰ǆ��ryv��:�£/�˻6��_�N�Y�t���I;��M�"�d��p~�5-��TF�g'�S�>�6�M��c��w�-��݇�������җ1��Ń���D'i�M�K�ӭ���>����-V�h!�K�� F�b�:��H�C�C)��T���n�Aq9�G�7�lQYC�ɱ&T�;)�& G-O*5���~9�P}N�V,��#�L���,ַ0��Sie/�ա�\1j�0��5[tj�$�5�.�[m��օ��JZ��Myv���X!+�Ky�L��V9:���Z
���_�5��ȔgF����XlxVHYEB    5fea    1830�����#Y`U��B�`�7��mPU��`��� �BN�ȅ"0ʂң?����],�swv�G)=��Q*
,yCW��Í[", �œ�AY�3x�8�C��iR�������긺���H?H��O�(���)x4o����9�0��C�#�<̈.؏y?�MAk+x�B���K�J	w���#vaБN�wf(�" ����͈Β�e�ʤ��q�K�I�$�k��Xp�@���)�B��}��m�7gm&����~z=x��������]�Iz0E�2d"�ʖiJ���7:�ƳIR���-e�}*�b��t���P��gQ��:G��M�Rß��QE�6�|3���(3dD������u��NL���	��fu�d=r)"���Ϟ���4I����P�?���	ܛ'�-`Q۔^�h�Y[�����������Zf�g���r�����p���B2�� �xz��ϙ�`��,FY0�d���_�'��g��0Oa��D�@���x�<8�����X�K�"�4�4�SK�?�2�}�;�����^+�`��H?Ls�mʚ�á�
��r�9ș�q.����SŭW��rcn��	��Ā1]`S�{V���Ќ��t�����ľ�#y�3�����w��Q���"Ӳ_�mG�0�����5�W��O5�i�N`-�-���D����ф=���Wb�w�ᙞ��6a�#�~�%�@�7)�S�����N���4��~$�u���^�v%�)!�q�~*GK�� '� ������$,_ՠ��f����`Yz%ʂ������zv������.���T?)�n=N��S+��Q ��J)��nm���%㲧z
0�/	��v��8�zl}�>GM,g�{���h��4��A̐�c��8�� �K��1@����9b����4ʘ`:�{�U'�;9�(;�s�����������1�͠���P]8�f���|�l�)E��Ke2#ˮ��O����\S��wܜi�`������IF�f���B��	�p�	fl	y�p��Anی�ҭ���p:�7�D�]�87H���+-�>G���d_��=�N�7��g;�.-t�|x+`+/ۀ�
׸�(��v���uw]3�0�l��A�A����[�и�L�$�7ǖ�:�Qw;�N� ҉ш<J/)�@B�T���>���Xi#�S�;�N�}(��)!f���)��zL�txt��1М�n�BQ�=���k0�	�o�9GE	^�����h� f�ir��Z�M����@�
������DnQns�|���]:I�R�@���@���2�79���jt # 9�H�Z�l�g�F��u$bg�{̺zs�|�E9��+&�T��$n�m���qT�R �+�������^��	FU�Օ�� 6���N!(�`�ZY�H^o�!����0��*c�x��;�FQ�u���N����)�K����'���K�;ľK�>���A�C"�y�C������-�e�������f��5�V��*%DL�y�����P�����	��+�E���NQ!�Ma��m�hE����Q�y0<X�?�|��X��%mt�h-�N�fT�����Kb<�y=�z����_O4/��J�#��vq���+�Pt߮�	Y'���S5��w]3��LB�����%�e�w[E�K82E�hk^�[�:�Xp���$�.�*Ԅ�6�5�;؅�J%j`����]��j�|�S$<3=}D4�.z�I���5�8����·�Ƹq}4��ME��b�2�k�Ì�
M;�Nh�#�V-EG/����&а�:�
�EsߗV����� St���I��%s�8���Q����b���kT��K�P˕�����7_wR�av)v�`@�:�����H�z��Ϥkg9ՠ>Ik���(���FZ�lh��UVN�^��Z5�=��\��O�_f)9��ܵf�{r~�������3'%�yN9���$�4�%}�;��W}o���7����8�Ԅ���iq�X*̔��uN��� I9ZP�e�cA�$ ���iw� Q"+:p��̉�8�A-�A���>�������չj��1�x�r���_`�J�A!��9��^�̓��Q�%�?�˫ m����Sb���]�}qF6�f���(�ev�LDKᢙ-��C	�L~����	S��*u��?xK�vEM"�\����2#?�1�a�%pl�<��l���u���?�_yeC ���k��/n�Q]o�Q�¶I}s{HG���U�k'o���.��%I�Fh�2b�F��}+�E�Ϲ1� ���a��k<��-��2���g�?25+�{�������ј��&ă���Z;�)�+���~�d�U�RTA�g*e�q�.Y��r�<C�uʠ)���_ͽ��cl:�ƈ�ջ�i�{+7%@&����L5�����=˰hl<�Uå��?O+�L*����r��%���r�ߩT7#qZp�,`��}�k]֎{1�&�[�Z�����P��{Ͳ�P��CG1#��r������$MN��a��7���D�`��p:O@g��eIn��t����T��U��PY�1D��Yt5M��:�Ri���{G��+N*Y��C�2j�@���ʺ�at���B ��1�V�=���e%�ϫEB���ͧ���t��`*���e:�ɏ�-�#6���!r�h��*���nl����\Mv{gf�'��sRFH�#,���"��A�z9��)'!���=��S�^���ݷ>�w�w:�u͇��\%���"�r��8φck�"�!^��2X��)ѫ��E�˺�I��i"=��ۀsu��b�wxg�נ��a�E���?s�2��m\���G�l��G'g�mE�t�Tv�i7���q�:BVX�
�W}�Z?�.�o�Ni�!Ÿ�>�,�@�PBw��ߺ�0�Q��,ϣcʭid�lL�W��l<���5:Uݟ�*|��w��,=��S�%=����w�4S�os�;����ۏ�>�#s���������z6���r�ܸ7	d�`�4N����D�G��mJ| |'��uM&���*��lXw�`f��Q�f��W��c��\Mm�9-�Tg^���2�+a\j����6��m�J�l3�g^"�=��^]��\����7,�&���MIYϹ�^'aHuTa^��Z{���E]�"/[�gDEy�f/2^>�6����{��6%���ƇV\_�u���2�.�N.]S��R�.22s�<�7]8He+�:�}c��[�.`�����bH�T���~qϰg�.����"�
l�+1'�v렜)ru����� ���ʚÆC�w�=Z�����\v�#�}���$$���1՘g�X�D��ؕ���N�0�[i6}���K�/}Qo�֭G/L�]�I�[ �>Vь(4Y�i��;���!��R-�Go.���z�	�#���8�r�m�hy�u�W��B.�Ġ*s"eE�����ϛ��(�Y���.w��m[�:S�
/��^���fڄ��iU%�!l�Ա���1z�wE��/Ѿ]��C4�
�3Q�4��w��ϡ�u�~4�3^��.h�0@�k!Nd��W���k4��L�,�YJu|�4���Ե���s�Oh5�6�l���ɭ�/`$!�(d��xX�n�x��/��К]P
x��`H^:��4�{U�hn}�[5L�/	�a�X}�A-�[΍:�W;�H]1gNN|��gE=s�9]G��p�`	�$�>�����"��}>�;czݝ��	�aY��k�R���SF����F�s��\r��p�۾����Y�$�+��?U�߻�a�H�~�3��,��W~�\C����l��6�x�%*�l�����A����;莋�VÊ�4c���:@mk4�B�"��ӝ2����C��1��t��;}J�����ȑ�F��(�[�/��߽� ��[5~�xjR>���3���rde�E�j���$�?��(��qc���j�h�9��J�!��J~�v,Ib�#l��c����-;[{�򕟘}��r�p��嫝(-=�R'*�\c�f��$�+�ynf�8��:|�1�v�c.G9-r�=B,���P�|T%��UO��7v�Y�~����N�QJ' ��c�\��S�z�[�߶��;1�I�P*��`�����dO���}Za�7����54�R�q8��[Z�5��GX�[��������S�����G%|�Zci�4��Z��Յ���,b�g}��^�ȩ�>�����TL�����<9(xZ����^z������u�[?�-&�B�,�$
��S�������&o��ͳ��Z��=PA��H�]ʘ�fx]�/�>y{3�	����G�y���#�(��"S�* �a�8��qg�ޘB�����s�.qy���vd�s�1:EI��n�̾��K���<M@*<�Y*���D��u�("2c+�HU.���������7N��G�-Y���BI|b�z'X'zO����NP��D���uLn�e�*|y�(՝-$�|���B�D.��ƫ���[4Lя����ެ����CI\�����z'6����� ��"��뜨�ب@�K�����e� 9�n؏���=�Z"�����ޥ���09Ţ@��9��p,�8�ͷ��%�:#w��S�b� �
���i�-�ِ��+&!��U��]?��J9S8��>�d��d���Uw҅���ʋ�H��'�2�Y��g��?�D�Y\��(עpӎ�� ���^x>����&̽=������I��l,I7�%@.�P�1�����C��F�˄\qƴ���z�����Ň�nԉU��z������0�nH!L��S���t�u�����,��̆��Nm�4�u��k�v�59I�5ЫnEl�e�yMA
��:�ڹ-L��;���VKqe�n�pn_�Q"�)Z�f'y�������A��8����E��3��[`g�v4��B`��/ټ7�9�0h"�Vظj�Pw��v=�m������e'�oτ��
X
z�J��:�p�6kj�=Pdg���Z�_��uV0B��*Gf�vs�c�NCC��.�Q�'� ��AbqF�҇�	.����DѦFn�4R����26�@�]=�H�+K����=�Fj��@�hTmKnD��yi�Co{��ؔ9baA��M��b�z�؟��\N����'��D�� '0h��_�;v�J�{<�H�=5Q	$�k�nTl��z^�y:Ƀ>)�&����."�[�ߦ`͟9Xl܃������!,���!��3�"r�\W{s����s����%��I���J�!Zy��LֿJ��ɩk%J��r�}�<�Jf��\.�܌̎�.��.W$Z\|�s�u�7WW2� ��5������pwmP`G�J�>��@���AD#�ַ?�X1I�L�1���X,���d��Ѯ-�'"����h�UPv�G��ĩ�d�E��й)�0x�}.]	���R�kg��wo��
ޫ�>����+�(�{���
�#f�T[���6�K�	��������/��}�1��`(�5"�IoFY�,09ĨƈL���^-L�Jj��|w�d�o��huT� /"t��U�E���+��Zۗ�}��& Hid9O�TB*�Y�n����DP��HϵJW�Tue}c��2��J</[ ��IT��0��=ÍM�����6�	m���)6Or{ύ�y��T�oє8����&t=�	�h��^����_e�e+���D7Lc��$��	 |uD����R����|"�ߟBE�GoL�x��а�������Mȫ�)�Z�>�*�����jW+n91�c��fp�"�GgDq�3�����qz�i�x�Ӹ���p�)����?�!@>�o��-"`Ԭ�~0H���-p�u][�G��=Ku5��Dp�w��V���"����qD��S��n��������K�l�=~g�$I��6�j�{7�%�ARY�dZ`���!2m��{�/� J{@B)7Ey��$p�G�~�����!�X�=7͚���"a:^Y�� ���"(��w<�*�<������R�Bŀi+��.J��&=.�|H'�M��?3��ԡ�`�t*��BB����X"rKᝯ��/�P�q�;l