XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���
�E��71�g�X?�?,��GWz�kG'�a�ߜ�c��ϋ�˲|�X��sN<��4��V��Jd���(�-�Ba�0�ed�˚�+�Vvk���Lz,�5(��u�,l�����ȴU�-F�žCy���R���޿;s@���܃G� K��:0��m��"�tЕ��B�����X���{�R�>{% ������e����ȍ�.z:ܨ����l�<\�e��'RwC�3c@� ��1��8��Kc��n|�����z�a)�L5�*��Y��7���%9��B��2\�h�����Ԅ�P���Tw`�)ֺy�_K�o�E���.s�yQ �)��"��F��w� �+R�"������!�}8��
����#'�4��~�m��o餲��^U%Cpk�ja�{j�2���]|v:�XO �gpQ��J M�V$}aI����X���f���j�=���;H�̦�m���X�M<�NNY�Ѱ��z,�]Ix���@CW����{�G�r)���p`�!-���(�~�\,��FP�V��43?��	S߰��!Á ��<v��gզ�s��fl��Qz�[�i�؝���d���e�S���2�%��Ⱦ/M�a��U��'u�甿�D��9d���#9w�=p��Ax��i�� �c�sF��Ư6��b
}�:�u��rӫo[M���͘�L|O��D����5�:����|Kg=WO=R�v�&�`	��vP����$>^�\��U*���Du�|�sXlxVHYEB    13ba     770���fFP�H�M0=� �¡Ч��� ��HG����p#�h�$�]�R�md�����5��R�1h酘V�L�D(�	�֭��S��D3�N���n����(:<�i���&-!�L�0}�ഫJ���f~��l ���G�D�q�[�W�Z�aw�3�C*�}JW ;��i�'�R{sY��t�ܧzۛ��"�\�q;�v���<s	��f�/]R�7ĩ��^��~淑��V���i�f�����a1�=� C�f��[щ#��J>J�'as�_�5�W1�K*�?�
��ǑJ���Vl&&֤�f����,,�����e!��� d�{Lۮ�_��:=� G=�W�߀���f
W�)��8&:C��2���Ap�`�j5��\ي������n{՝���%V5�������?��r�.%W�!3��i��MEI"U�<�D����B��԰��ʜ|>�[�;�Y�u\�KlԮ�0V��:Q��)
"W+0#�)[���r�)��'���#w�[?�%a�f��J�E*�r�U���R��,L�3���Y����z�
�ʤe[[��]l�~�����m�/���b��O��= lv��2�#}e��Qb�6kB���h�(�#�b���u_2���&~�|���8I�ǎ*�C�ID�8D�>�D*b$���  �Ƽ5�P��q4K�h��X���֟�I�~<�I�i7w�6����eJ?��?�HR��6��=�����B���!΢�[�&[��b�Į����� ��i�w��Z?����U�n�g����-�ow�g��A|ڔ���Mu��������l`�M�d������t�7�ݬg�Ѳ�����ǭ+<��Z��QJI�~�v;�z���ܩ(��@������g��q���Ǣ�<�]aj �Wb�K�+�/�����),��vꏟ2��wm���0l�� ������D�r^'�2���3�vES�d�V^�Ŧ�5#�-@���uT�5w}X�E�dA`X3m��HC�x͈�b���3��:=�+	����f��#�\(�u� ��k��0��X�$�(<[e�뜓���6�GzPf��!r��'�F�-��w�51�~1 �{8 ,f�n`���r��^�L|V詿,j���ɿGo��JiZ��ñ6��A�^�|!s��J�<�5�E�м]ڽ|OH�K5?K������:q獎���P*r^��(<�=�H�4�g��ТP*�W#Z��j�(���q?%�j���>-�n�F��u���.��&�Ϗ�Aβ^o��{�i��:��У����X���($���T���"�O�@ w[T-2ƌ�~�¥��u��~v�P0���O�5<�Ṍ��VI��hH�#u���iQv1�g��u잯��2�Sƒ��ČR{γ]O�%�ɫ"�H�z9=zg8�7� ��'��P>Y)�4?��=?6z8g�k�#�n{�B����Gǥ��yc0N��7f,}�p<��=d���PF4�Es0n���X��\_���#Č-����|OJ*@:)!Mعn��Cj��Nn�Lq9��"K��Rd��k+u�$l��T�c�\(4�����k��1dv�%w@��G�U��]3�~���{�Cߧ�9�ns�����'u�ș�K<�e,#͸ܹo2��/;�e����u
~x�K{��!KKZe"�����cF�$ "��rR�E����evJ��'=p��͜��H�o?1�����[t'?*E��`>�@��g$��R�R�[�y�N�>�����^f��T�ώ�y�����[l#���(����Z�Wl��t��U�\Ʊ��E
����� O=%��J��6�*BG����X��I�CL���[���Y��