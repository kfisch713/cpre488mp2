XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}$ީw�����0����o��u�	��(T�[u��ȑ�^;e0��*ǿh��?������g5��7�pj��N�l���G���@0s��#�#�pzd�
_@����S7Ţy�?��_�-��1d|2����1rd�$��O� O�8�j���Nb����������L�D�� F�.K�E DV<��. �����C�d= �g�NѶ���-A�=�Ո���9�jv�� ���,��- �)��(��܁�li[C���l�X�]�Lt�xU��ߤ�w�[w�v
!8yy?�~���~�h2X���E�0�H��T���(٬�G��`��gY�]�
D?�K���m��!�z�Cr���W�v�_7�ق"*�pN6k�j��L�x	ꕍ׻E{��+~r���M��)I*Ӿ*ɚ^����db�r8��O����|HXkx�r-���2�y�>���$>iu>���
KЌ�!KeR#��̍���Ub�ѫ��8 *P��O�4���Y#��Z��Ro�` �>$.\ 8f�12�G������41 4|�B��v�j#��F�p�_&b��xi��
8�ZE9��f�
�O_ڪ�+��-�р�"��\ M�D�p\7Ѡ�g� M*��^�e3���k�b���I�����yi�Boq�>�.`���*���]je/�f>�)�ٳ|���/�/%�g��r��Z�c��x_�T��}��*�~�G(8Y�f�$�% �N���?�"�2�_땁,�5�A5��h�B!XlxVHYEB    1959     920~�ڑ}��d�nQ�>d������P��#�k�<�<t5�㼑�Rd� �f�I�k� ^����E�2���Y�,R}�NU?����SY���'�~�zŋ�8}6�,��(�3��h��J-�øV4��RN"1�d��� i��L�E�X��Ǩ�#7Q�q�h5����._B�?��4�7�~�,"�>כl��\]��%*|�)�W;�������Xd�C�c���_�s��Ӥ���$,(޼G�����7d���t�]W������IT�W=m��,��vk�H�x(��`Vy/ac����Y��_�����L"��_؈i��.��f����v�t8:J}�^�>�֍ Y��`������G嗥q���hZ~H:O~n�V��5�)��us��B�ކE�Z�����.؎k$� @L����]�>�bh�L�t�@��ɋ��Ngun�WK	��-
ͥ&��Ŭ��b�~f�'�2�Wt�K-�wp�c�~��)�G��U��aE/�.x�R@.��Z�62j3[`��9��R�r���4���]U'Lĭ�ѫ,������'Q:(��}lP<�2Nl��k�r��LT*�=[�WA�J��
�b���'�v��Q�o.�_8��2�viҿ�X�0K�el�(�����p>�
@�a�������y�8R�����R��ā�IAK���u�B�"��;����\09�R�LIU�{D��8�׀�Z�t':��"t���|�����7S��,�E_T�77���h����2ۏO"�gs����06;����j��2k�D�Oy�O6��@~��;����C���k��T�x��w�CT��i�t�Ź���UA����&!��cq�WM��5L�����2Xy�WmJA~�$T���v��y����BD�[T[�o)&୦ʰ���rxu���-�t����_?���r����J�=�~k��,R�k!<D� �>x�/1���)�����B�����K1vm+�ԑ��3:l䩎?�3K��q���>AX-/�I����������Y<�H[���GxX�ƈ{XIq� W��ր*5��o�*Y f�)�y(���>�6���ɗ���SVJ��)Ac��uaW� 7r&��=�E4���/Y��%�,]91�y-3)C�_��xR��_�v�
U`�]���>a���n�HY>�/la���5�N��Qɲ�Da�9^k
h�f���D�|�L^ˠ�4GJ�H��܇_��#U�_���'	�Eb�hr�NRb�E�\x�B���������u������rA�� �O��&�M���_9���C"ү!$M�_�2PtK�"�$��kO�ۉdl�����M�Le�d�%��P'�gæ�ݤ�N����aX���p���p�7��"�d�ݬ,�\��l��
:�w�d�A�7���#�Y%OK��5�j��G�Ni�@�`���Wi�K��2y0�4=��oM�#'O�t(��r�O��䩞A�Ù�T=F����bX�{Ɨz|(D9hqLk���)�
��XEn묊�Ik�d[1�YC�o�|S�cr)�|��"KN�tۺ�"��2�>j�PPhe����qA:�b��O�/�����g��<�dQ����,�x~N?����e��O��qW�!��no�P���+M�1���7�J��%������`GG��⬊ltvB��L�����!�={�P��}�L�_�Z��@z�@�Y��M�	�_'mW�~�?{��ֽ"����[N�a\m\��,��Q GM��,�j��9���HJw��vI-��B$A����U����g��t��k�J�{Z�7���c��Y�I*��d<�$�i��پ���O� �>۰]�I`�F�Qon2S\���n�1�R����H
� ��U�r9���4Xd��t�k$�f�e����пUT�k�;�>oD���u��$Pg{O��5���lL�+}�<��YY�,nֻCKS��[�R�gg�\ �R�� $*���&�O"nz�c#R�V��ͫ�H�*p���U%�1K����E�E&�6�:�/�a��=�7~4T��f��ƀ�p 2c(��ǎj5OĖ
�-����#��wԅ����B�(U9S~�� �@��j�D~w����}���8��������d��8�Gk=���)�U�8�����^����0����V�6�u ��Ța&�/��f�c�4�QG'���yp�i�m� a_��(�c*L�x�������7-+��q�����BuJ
���.�?8���Ɓ5,�M�^�l$�