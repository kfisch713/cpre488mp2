XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+���05&�!�i	�t/ B�6��:a 8fTJJ�Қ�'�wm`FDŁ=�H	:0�.b�T�w[�09@RH��Q0�s��+��4yP3���$=����rgo�&��WmWEN}��As-�F����a��Z���D����j�#��D��y���\��-G"sц�S���-�5?N�wH�f?��$ 2m2`戗��ڦ�y�Ĥ-�k�MD{ŏy74���=ܮ��D-s����a�o�����
|�2�vh	��'��t�4�&L�!�q���b��o2l����V�z�87�vQ����vn���t�i ��*�VwN&ވ��T�?��X5�yK7$-E\82���@U��Q��/�ITh�s.�d0�PP����U-Vx�� �6�ì�M���ӄdL���h^��y<�K�P]��Kڤ��*j1� ��SZ��(4
s�Uy�h�5007[��T�|�t$��I�����82�XM�9����e�g�1�;H4:6��4���f�u�c�͕�Q���G�VQG�Nk����Jba5�����r�e%0�f
���(kNL�dQ�	�vU�e�ѿ�eD�8�n`��B<�$3%�}2�Z�P��h7^��\�<�Pw���*��mL��$O���y���ҹҵ��(�YiB��g^ai}��'G���2��+M;�Q>��|y�J��́mXa#XOA��/8}o�K�C8�+��p�"^>]vx������ė>�/�I���.g9Fa�y*T;u�>��c_���9i}�%5`�XlxVHYEB    13ba     770W�O��Y�<��^�{��wC�9չ�3Ha�L����TV��U#(��h�#�AߛEWt�w��K���W'������-ꃚO�ڋ?A(�UZ+)���0�BZf�Ħkw<vަ6��4����5Gfn���3��Ͼ��������qQ��_�#��̦���f����bA�������Ex���j���������ր>�`(4��ȯ���1w��i;���G��kr��ˎ��lU��0雟��]�#1���Q�8j	��y�i3X�f�f�~pϫ�sܮ��e����(IZ��'ge6s�UƕU/�2 V[�bY�R��4#w`�̈́���i<�Ҭ���`����@��r���&EJP���A�� ����?�׍�P"i�Ǒ�HÀ�d$�|��QF�wz��f�-��M�\kZf��#n��sdR��m��BE��N�#/��z��^�{±V 8�$�`���l�Z����ݙ�� ��@gB�cS�Z���8�ܼT20T)����
-r#(1�� ��]8�=B��~�@T�Jr�f9Ŵ)��n�� [k:��$TG| �u�$�}0⪽��m�c+� �i/do��H���\A����u��p���?���A;�'�Mg�6�0��
n����-lS�U����0�[_��/�O~s�A���D�{`B6����Zb;I�pE��
ڛ�/��Uر7k��A`�1�Uޏ$�g��Lv���?_V#�U����h0�� ���*iX��.�"��o��#!;T1���e�`I��s?jA��Ó�;o~V	뵹�:����-�t�_v$h8�I2�z,��Oi3=d8�ȡ�U��׏�
�U�ј��5�oa����u�IBS'���oIn���	�f�~%y��e�A`;P�)��|����ҊЭd��&�9��*t�6fk"�F�O��^|b��	��ݍ�֜���r`�Hm.��ړ�
ň�`�qr��C�=��X_�k��� �2BYj��Q�0;���A���p�t�����X����^�@�Q��;m��`�C��#c*3����<���{{6��^
���Չ3m~��|]��OGF�|�Y��r��� ��E�H� ��!5Hyi� �7��`?� 	�"�FW!����I�i��{�8m����#\4������X��T��*��K$�l���U�L���H�Rr�����X
"���%�D	B�n��筈����'��:dҨcR�Ҁ_��+����ܪY��_"I�b"�d�7j�0�׏�=�L���x���?��|���R�.�Ι�n1)Ք ��90��]Hr�2@���;��'�|�`�ʶ�;��y��d<q�����,�k�A"����:j3f|���s�#��(�x�+���D��NUˆ׽���r��qˇ�>�8K�gm���j!H��<�S�\�4�G�[.d����5S�s'�]�ՙ;�C��%u,�Y��c�������e�kA��j�(p�6r���Sz)�z���[�d5����=aGZYB���_>��������u-��rތ���/"�#Fta�7���o���z�v<|ß댏��AQs,ge/��D'��A
�h&���`}�]Q�8�Q� <U����F�	9x���ۢI����b!�Q��z���;h�0�Q�P��;@��M�'[o`��Il�K�����Tn����8A�K��92��?���S�j;�1��z5���50m�>�2��~jgtS�Z�S]*`��I����L^j���ߏ�p]xa���m
^���5�BE�Ă'] rULb�R>���8�''^�mn��Y��$��� i�e�,Ќ�t��P�:c��9�����@��"Xn�$��Ҿg��|