XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�6�7�ڻ���ŗ�c����ܵ��iƬ����M6;��f����`�vJ�[-x$m�V��ǩ�n�����mE��:X��4��5 k��u�ƭ7�Sݫ
��B	���d�x N>-�c�e�ӊg_6蜳�(/M�,稥J��̎�X�p��A��[f�8>\�,�n_�8q�l���f&�D��)�fJ=_Q/��?0N�6.Di��;/+B`+2༘�Gt�=�O~�[�pxq@�Y�;����N0����c���]�'b��[L�J�h����ZNN���MniTS��ɒl�����s+��(z5�\�2�;}�]Iŗ�(k��}!�
�~+U�qz���En���(F�GF�ۃ�܋�kO�TgyT'.��/\��Z��Q�A��ҍ�ˍޖQ��Ĭ��,��Z�q����S+;�[��mG1��RY.��0F�9�`���g������#�����³tH~ϭ������0x�j�7�jT~�e�7������X��-R'�Ze9�JĊ�kR��B��eBc��⠘�����j�JL�f8;��QB�9������ґs���9��t%W��ku���E���Μf�M�d7��`MU��?;��q%�Fk���˓P:�E@��%]�����z]Fg�_G�G��ô@�:���b0+�iu��r�N��?��4��(`�S��CBX�<���x�k@	�o�FJ3��~�?�2#5H�Z�V�r,9�h�MD0���4O���4~�nJXlxVHYEB    4284    1110g-`?j�6��-�:��q{�h�3\]�*���'��������nu��`��]�6mL��`^׶��="��{�5ʻ�r�,*x�G/�@})�`"ɻ���������}7�+Ř�L�#�iD��x�'�E�����Ci݇w#kVxGS�/���tN��9�����-�K:�U�Y�ߒ�\��/6,��M�(H;��<|-�6�+Шt켔��E�AF':T"�z��nB�ð�\���=�q"f�5Ӎ��v��p��,F'0k�FJ�>؂j�j��YXØd��2���$4�T�׌z�0P��Gv��4��[�/�,�NϏ��M�V���T�A�n��D���Y9GBA�1��}"d|I잍�-6���@�OKΈRƙ�3'=�c�XD��ǨO�3��j3�&ȵ $�����\�KcqXj2.�^V=N��f5LeVm�ƾR��b����7�ĺWE&�1�߀"�<^mt�s��+�,��b2���-����÷���)}v�s��KRi>�\yVt�*��b85��}bX{���/~"O��-#��'�����ҫ�4���z��8͂��ߟ���
���R��`�q�h�Rs���A�Wb�2b��6s��][mn�I�ڿO�A[�3��o�!*�B:��G�QQ3�5e��w[�XVCl�������e���@��X�����ef��WD?U&_V�7y�,����RHNi�_ą��QfG0�Jrj�	Hۺ�aR{%@ڏ���<�J�Cb��݌�B+'�%�)�(@,�h�ß��9#Pc��h���d�E�_�ٱ�K!�4��8�,J,���u��\1�Zܓth�L���CΣ1�y
'NZ�8=�h�}��Ř)#�m>3��g^&H��ƚh�?�!>s6���@>�G��Y��|n�v�_e�$hi�����ӕl�i"��Xj��w�9d��6���J���H��W˶iH��-ڱ3��X����9�M$�j��{��%a������I�hp�����⧯x�Pn��B�P�D�W�lܴؕ�*>����CY������.�(e �w�8��X��KTs�j��
Y�ղW�~�S������'C�IK����,i�jm)V��=?r���$ݣ�q�?M��,&�B7�r��υy&����>{�:�DW�?�U�ɏ�_-�Q0㺄e���Q53Ln��h�-���'@4��.I�����'\�b�b��2�O`���S<�] �D)��1�'�٣�������3�ѐ��,_%�q8��9��Pd�#�`j�ݦ�Af���f��	?٩�8S�"��f$�h��j��>���V٦��
�)�Yp�tnZ��=n�R!{�0{0F��k��J��ޖ�®ʯ+uTw�h���(s��)Z4�R�c7����=1����(H�,�;��̀t�zޥ��ul�g՚�>C��BA~���fH�IɿC�
1���z��Y�/m��Ե�=�7�4��N͎����`�'�Q#P�7�C��,��NG��4��>���J���oKʰ<B���w�+y�y�#K�Q����\ag�
J��yQv�^�	X������_�o��B�Id�����B#Ea[��M��(? ��A��1]�*�-nE40Ĭ�ڜ|��Wt�����U�c��{p����h�Ḩ�:����>� ��43�/�28��w�Z���^HW���n/�=|%���/K�8���~.E����2j�&���h�4=t�j�Z�!虪?�6s8go�� �DomC���X��b�r����
o\�y���t���Hi����R�se�`7��N���� �0ZQ��0�Gܦ�G�M�dV�H�����M|�I�T���G
��ې�l�Ď���")���Ih�1�.Z��ݢzM/��V��P���.@͂ί�߈[����wS��o<�� a����pͳ��f_%q��b��i&����-��*�3ͅ��^��I�2Jf�B|��q-��Ҋ>�Y�6�3��և��<�$N�43��]�C�7�.G�Iꁾ2f����y�x�U 7d�|p9Sy��Z�S�Lu7z��d@����B��c-�UD�C�=���N⁄��:�nu���Nſ��z����D^��2��ax���葓���%ha��K��2Q�@���j4/Xa��m&q{|[�.b�"�;�l�x������%²@z]T.i�Wpf��I	/qۉt�ZeBj�=ra�"��{ʞh�P�.�nyP�^*E4r@�N?�i�)�A��뒘��K���"��_..TQ颿�6��[�7؞IC�����Q�+�ɰ[���$�[�@�*Cl��弡!'TذL� B�C�ۀ��P�����$g޽�0�T��I�=
�3LG�ue�����m�ƫS�^R.��%��(9�&��2�C�;ey�ƣ;{���J��f��9��I@1q��tk.#�񖕔�_H�&
��U���Ey5ޙ�"�27s���m�<��(�����9
���Ec.��M��.�n)�h�8=�P3�bG���Q�?�p1�F� ���c�v��_���@����^�>�[�{�8+��t_&Һ���an��V^��s��`���R�Bh�g�w����������U�?e�u�mQ�?N�Z�d�Y�-�hQY�qi)���ڣy����f^�w��.�B9�C̃�����\雹��S�M�~w�l]�9M����C��F�ulM���wW3�y1*��k��A��A���T)��9��1��أ~u ܆P~�J8�:8@����Q�F�Xq���z����h���؄��g�<N�f�K�+Mߜ,_�����.���j�A�b�їKj��r�k@��a! ���]����q�Ǝ��Ϯ��h�&�1C�8j�4�f��\1��Di�yI�P�
]�<P�xK�*qHB���|�Cy���$>_I>�5�s�*�@�׭)dyǍ k����)�FiU���m�y�,u��J���c��b����jluK`=I��R�tz:_.��ZƂw=C�AP���� ��,S"}.?� �|2$���8�M�
j� �(���;0�ٙ�?ã������u0LH��������W���$��>F���sB�V�>ǣC�HU�Vi�&e@��	9�~��e��j�ZRv�dEm��keV�W�R��X�G�OU9}?Q�ѳ��DK�%���%Q�&ҷ}�U���aa~��X�xѭP�6B��a*.�A�F6x[qh�&�_�q���]�WD_EO#�AO�r?V�G'�������lSC�pR�Y����h�}�h�^$G�6�'.��}v�4����H�%X�h{i�o
�Tݝ�����C�MfQ&do�r!km(�2���u͘��
�|�X�¿f�unh#���1|�'2���,�uU�@�2N֝�fE�����D��x�$����ۏϷ�1&҂�m�šfy��3�������'�*~o>���sʵ�h��n� ��ֻ�w*��=��:Cr���K��)�w��9�v��;qbP5�����Ъ��v��٭M��R�]�"�����3)1�b;�L�������_+Qlp�
�)aڑ,�g�gÂ�ι�X]�F��@��O�A��������|���
��j[�wGŴb��~��iyJ���� �H��RG1�G�MGb��3�8��8q����\w�Q�#�q�Yj���&Z�8��sl6è~jy+A��/���AYz:5��#I������8(r�4H����	)�G�F]?6(�ZI��h�|#� ����w�S��w��N�-�em���M�u�x���z�ب0i9pc��DzM˘]�j��l�^�U��_X ���.q��|"aE�˟8�U�/G�ȧ�Tm7=7FS����#TS����QT��g�Փ��D�6�85h-u&8[�բ-��t܍}A�����d}���5Z+oG~���`���9��5綞�Ť+bNf��L]��H4�GhKi@��"�R��Y�Q����؁�;*AR�]�m�3�S7oŨ�Bh��A�F��9^�f(���6إ�|��#���>o��B�dxñ����8�~ԏ��r�gO�Ӣ�^5̚��f�N���:]1�1��)^_E��̓n�i8%�C�Ġ����\�o�m;N�� 7T���v���:3�����|H��@�W�,����%� �U�9�y<�y�/_vᎁ̱ ����Ŀ���ܾ�z�]�ð�謣�X���~�O�&��A�w���7Şj5��,��$\���J�G��O�א��8rk������7���_�-lUdi�n��C/32��v��?x�#8�3