XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��h������D��Y �]w����t���x$k�����f����%��#�1d���aC*`֋2ST.^?@�����+5%�{��AV��/�;>|�f_
�RP;*qT�X��t�I.�I��E�4�l�M5��@��9���$�?p�{uH{�U8����^V�N��0o��=�>M0���ٓ*���4Jǆkma����G�����+�5��E�m@��c���"�`k�[��[�몟�����ة�l�p�.�]}~F�����`�n�V���M�ˠ~��X���S���)�@�f=ԟH��. X��	&�kNF^����`��\�r��Ɗ7���	 ��#,_kvm�9�L�"	�k�,�8,GQ }��R\E6WR;Dzq��{  �dt��Z������#E�e<;�+��yzϩ�p/YR�Y��ڟ�%�r{���\��B����z�*����t��j��.����C��j���dUE��;�Ҿ5��Լ^�;b�6s �zmG���թ�Z {����/ ��5w�����_{��p�l��+���M6�ک)���hR�%��R���ra2���1�a�0:x_;�D2���T_�vVw`\ojYL��לl������3�];24��XsAd �'�1�> �rjy�JF�bTH��c%�����;aw��~Z�j/^�I��}���P�8�ꎶ�In�0\ �oB$����2*�N`L"Iw���&7��ut��5�R���,1XlxVHYEB    1421     7a0:Om_���έ�6����g��c�#Qs�ل��ƍդ���By�A�g�s�F�`�KfX���b��=^�^�`h��� RF٫W[x#�f�1~�8��H	++fs_��;S>��@�ZM>�{ש���8Eu�bj�Q�8S��	]�, ����fɚ�\�ꋫҕ��V_N������
��^�M��X$�U$(��j`�&%�G�Ţu�n���$ˤ#���2���S�=�SG	�i�Up��yՉv��ǯk�.���$�aB�\��ez�^�h����B��4���҃O�-=�`��+�wz��3���r����B	WQ(��0'
Ϊ��!GL:��U��4��sC����GC��u��W*V�\͟N���I>.��@����o|�.K}4�`���:�����%qn�*ص���2鯅n�,ɯyB�!�X6V���Jn��0���<�V��թ���ӎ�r=!��.U&�?�ط����>+y���� ��P�Ȼ���0[s�f����+��M@���߸q�=�)A5�`i�U�	�����+�d�#��H#���`n!�e(̆���]2#!kך���,�&SL:0�����9�K׵N�	���41��]���_ĉnl��( ��+(�����p� siȸH��8�����O��R���:<�Q�V!�s���R��م�u-.b�RC�'��A\@g<K�#$�Skx����c���=`A��ؤ�I�5��`0�~�Ձ���SS�%��(�#��Lu	/`Y����-h��R�����8V��4�H���<��'J��0�GO�u�(Pf2q]ĝKn�ū_�A69��H����
�~CG�_�!��2���D��� ��R`74B�l�{�lg�o]o 𱞈H�d, XШIi�ԃ�S*\�p�t�l*��U�L��O�B{TX;��|�mX�r�d*ۖ?����2�m������k1LղϽ�v�U��Dq����DoKۄ(Cټ�8�
k[��������m%�<�2�eDU��q]>e.��E�(>(���ʈ��B����	7���������8z�(l9�`h��� n�ҷ�2m2ɔh>��\����T(Ű�c�+�j@�(z����A�LyE��v;���iQ��(�Uwk�(w;�^����{���i�``~p��!<���{�^:A:fhu<���[����v,'l�	6nx@���q�8�I��gĳ���y���E�x0��:prl8 ���})eP�_���Y�wƈ�{��F�5�'����e���GyzS�<��0�`����H�*|�YHj�Sτ�?ߵ���X�-T��߃��j&l�Q��0[�Xؖ$.��>�ˆv*Q�/�L�crcZ�v�[Ȁ�(�s(\�L���z��-l$�	����~L�I�j ��U��bx�W�K#�U��Ao�O�d��xI<����=;{�E�<�C��yf�� ]<=Bm��o:B��Ϛ<���a�q�6�ߔ'�JS�x�F�j���X�eLݿ<4)D��odD�d�k_�PY�Up֮eU��Mv���=����6��^%P�s����hL��S�QU�+��|��r���>�}+���Y&
�
x�� *G��
s�22p�۽U�QsA�O@���w.R+�tP^����%���	��T�|\��>)?=W�y%�]D)�!,2A�D�(��>#����ȏ9d�3���:չ�f��t� ����"��	Z�����wϿ�o�K$�6����b��2��9[$il%K��L�뉞����G=o���Ȣ3���j��u4���𝄌��x��$CM#��Y�{ͣ��Lc>�{���a�w,^�`���9�Ѫ	��|>r��j^�*�����g-bwq�g�y�&KS�nRW���ߎ���G�6��$��Q*��� w!'Zs?�8��Oƥ�j�