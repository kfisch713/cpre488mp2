XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v���ۏE�N59U�|�i�b3��'Ӱ
�Q�/9ڗ�P:hߐ{P͈�+m�}�N��H�"?J5���j.�x�m�]i�ڇ��b6���������5R���b����z!��<��ɇ�<�b��V�8[0#�G�'�J2�+|����v ]����I��-Q٬�
-�|�B�.����h������,��E�W�_���Qge�EA������P;d&'��PH&�͡���|`G	i�"�oz����ߑ��3��q�].9�9w���т�J�;�"���f�������+Iy��ȳ�W����?��^'_�r���3a��H=W��Yskرh���I J�8����0r$
�5W񝲛����_#u���sl��A�L�h��i�	�J��Z��}v=�/�϶� N���C=
r5w�[�ߝ=�K?{�f>�X��e��'��aV��xpp"� q��`r�A�T�9b��^��ds˙�_nn�e�u�s�QuW�)���{�ේ�dq������2fM��bܝ�:{�,�s���R�;漹w�}�Q�����n(��	����]�q�}$�� 
���_O9�NT��4��1�U7�I������d�Eb3P��;gd�J
`��1���[œ��;o����FBI����^�D�+�cG�n�\;�B�p���N\)O�3Pfʹ���~�#G3�:���܂E���5�mZ�_�n�l�}�#�jN=�������3N`�#�:��@����M/�
��I�.>�L�JXlxVHYEB    1847     900�Z �_�]OwfU�Q�Kx��]{� cxգH(��*�n�y ҝ=���:�: �	��A#��O����,=�#.��'!X��y<���%0FR����W�Qg�H��.w�e�Ae�b��[��^v��sy밽�(Q
��\#�W�o�@v`]�̮f���=$>�!
@7������U���S�2f� ,}<�v+��r�#�h� #�d論&��HI�Gjn6ćM�,6`}�eM z���Bh�&I���� }����[uͶ�@HW���;����K�� �i���J�-7��L�(.?���i��}isW���T��s)+�[x5�Q�4�ѝV��M�`w�?d3(|́B(���Cv�2�"f���2�¡)� p���pz���(��}D�k��M1��5!��#3
�����Ձi2f�xDyL�\Ы��G�s������w��d�<uz���>��9�B������|��v�����)�_O��3hEC�cS+�Ӳ���rH<5'j:nP��f��,^�о	j��e��X��� jɹHE����Q]�?:=���ق��)��a�*^p�l�(��=Z��g�J���
����|lڣ�8��J��x�ެ[�FB��0�07��1�0YBL0Yӣ�@㺯&7��Ҥ��bQ?��i
�v3s����n���i��B��(5����n͊S�:~�ܲ���)+�o�?n�:�?�O~@R}{4��c �����C�eu6)��&C��Lwә�r;� aX�����q��.ӿG�8(�zA C��s4Qʖ��Fq6�a&m�&��!r�bc-�Ǯ�xy���&����k�t�[��[�l1%ء�cR��ك�Q��D��:�a����&�$�BK�3`:�2.��F��	ݔ��K�#g��П��!���*�^JE`-T �c�p���+�[�������\%�W4t����|ǚ�u�'�=ӵ�uQ��曡2�VK�|��b��kՈ����),���7��b}�����sP/�6&�㕁]�Ou���q���I��0�;�@s����8^e��\ׯL�,z�祖�t<�0b�t�4I��M7Z���O�w�q��p���F-z��-�K�m��3��mgV�\��T��Foqn���*�ۧ�kd�����e4�;p4���4��c�[t��+�T�}$,�������6~�D�������N�NY�k��$�u?F7�sK���m���Npd*������m���z?���D
e�Xգ�_�{ź��I�\�hɯ3o7F����+�J��KH��:u������ o�Zx����B 6o�`�e�0���o�`�s�>�$%W.th`��՗�Ij���*V宗�g��+�q�ր�ԎUԹ}�?���/���GGx7kJ�N�6��@j�[nc~}q��C�?�\�.�9@��e�ܰ����6�r!M«Ouא@�}9ox�L��4u��V��a��w�3t��,2ӡ�� m���p��HHP�}6R�*�^7Z��;GU���X�9&�)�^���Y"�J���1�]���g��H�<qi�s��e��jW"����;�N�a��Q�Q\����D��2j]O���=S�@6!��LU7,e$X���I��:�H�=��䘌eye
��}~7���[xNP�=�*Xe�=�'7+�3��
���綨W�z��;�C��+n��Z+��<���:��ƾ-�������/�@7�h��?��[)�7)����t�Ee+��z�U�xl��|?��۵=t�?]qL����B���k�u@2�A%)b
��.Z4�Qby5�����Ʒ�*�)���G�_}]��!�93�z��1#�Va�c���=��X���l+i_�e/1�q*.�bQ���,R�{���vC9��3ek<�2���jF�i��@+2[�)؈q�V�*�̍��酡B92^�a�t���t�NJX� �ǽjj�=4Fo�>D�'c�P2Z�c`�N>@I�osM0���B*�q�qn�7�%=u�V�J�☓Hϵ�8H9����:�b��j��p�0IPƦ�+A^��7�C�WUw���`�M甋V]�H��7>nS�ǩE�}QN6|�O: �9��U�@1���^�� �X~�KH���e�O�U�[�8��F9.�t�I~+�6R�`�ʣm/T����E��_ �9@R|���H��i�"a�r$�U��'�qĠ����vl��de�I�"c������%���ن�������{�g���Y�����