XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���f����ub|:������ǫ�s����<�������l��D��� �v*S���x�&�7'�n����\�S�9xRP}2૚q��d�0�@
F��p���Px�v���j�3��ҋ ��U��!L'���;�'!1i<���7R�\dɔ�`LM�?��K6��ri�[�W�Ys��x��$R;��/����W�pTc��a���OB���IbV�2��*��pQ@#����L�?(�oF�7�9[�
�[Q�\ZW}P�X�n�b/��+�WV���|4�i�F�Qo�m^�A�;�\+�ہ٨cA@���F(�\ф�8�JI�l-U�_
�Z澍U���l���e��&�K�/@�;����ir%d�)�b�{(�0ŷ�7k��f����$v2I ��~n�6k�\	����5BI��8�����3��M漸C���Pv0�u��Wc�v�XD"�h���U,@�����ʖ<�r8"X�2��K�j/�y���#�z*���K�P	����[l*�Sò�E������Q�^L��w<75{�ׯƾ��a�o����F� g�-�.�r����B� �09���G1��n���7�1����`P����X�n믈�V��LI�$sN�� c�$(V��<HE�Z׻5�@���0�+������mczAFFӟ���̺<B��o�ڋ��!Q�,�8�R�-�~�h�Ris�C/yM���"��7��s���"B���F����&����$�����аy}�p�w��oG�XlxVHYEB    5224    1740B�<f�*pJ�L�uj��ϋdj�"T���-,�ҤV0}W����D��K�/9�F.�"!���&Cu	�b�f.7I�H-Thiq>2*��K�Ǭ�A��zR�fmk��Y���+C-�;R����%˜v��)>M�Ml�Ϗ�p��`��]����"��)�v����5[�A�X��冖-�(��5�[N� Zf�w�5��;=O"�D��TTڂ�Ɍ�H���+1�@M@N���w��V����
F�Y$-�J�C�H��9�Y�_�.V��S�����qey�7L���׷k;�����(�5�����o�)���2���(��^��C��E��k��,ۅ}8��?#V�) Lh����i~��	��Ar	AciϜ��&j��1{�*�w� V��>��>�x��\9*Q#�,F��
�bMf&�p�X�-�UЪXF�+�m��Ձ� &!n�W7~�?>�zd�'|��b�J�鯥��){�b��8���z��fC���="9�E�)@\�v��2�@��:R+5�Lä�	Pe�n�sL��f��d}�XiZ`,�M ���������c�[5��7(�@�ɤ��ϫ5E���-]�S�z	�'N93L�������/%���*X�q�,���M�Ŋ�kԭݼ�(�V)�ԛӔ)��t3��S>�%�����C��q�1�X�-�O������!�\&j� ^��u5"�'D-����װʑi��Y���	�����cԊ�?;�446�yŗ��.P�4���16�����
��C@�ͭ>=Ǜ��g�k(]�Ǎ��qd	^b�z�Gr�T����������m��`5�/�V:�-�Ջ(oT.�ۛ`���p���lAE*�t#@y2�= �z,Z��r���y�8R��;�%��V���&�����8�R,�*W�K������ xh4a�]��L��b��iЁ>��t�l}�@{0���rE#��O�)H�(��w���E/vVX�1�����wB{�@܅��N!�Nb��3����'��BOp(�#��Ȟ���m�U�u����S����V]�ҙU-%����0��U<�Ri���� 3��j�p\)�i�*Y�qҭզf�Z������F��X{.�����9����by��WY����f$<�_��Z�\Yn[����l��n���ɀ}��$���wSx�٦���� ^R��t�fZ�P� �i���4��W��`h��웤���H�mi��&�L�:be�$��U$.�L^��!�,�Hi�MH&���-�~����U;@C`j��&�?ԉS�7	E��,*Y�먤/"��Ɍ� hS��5���YT@ɿ�V��]����wFt,�#�����i1t�ni�4�cB�\~����q���8�w��M��b!g�E�֑_"�]�0�օ�e�x�y�`�i�J�;2�D�f$O}�I����d���'g��{���HzT�Xf�Cq���z^����s���H���;���լ���Ju���#�Q,���zB.$XK�e��tA���}푴�~N�ʵ��V~]Y�(�ȰKX�e~�����Z��#B`)��@��S�܍ֻBzW���QC��OE��9�5����T�j���Y�@�Q��K[Gh�g#�6�����=�iõ��oW��NoZה+�ұ���V��� ɤ�
�rP�#�WE87^b��#���B&��
�i�Ç�T���p���m<Y�Cv���y!�����lHM�1�e��G�T��72��S|�PXzʍA
u�b�w�[9 �6��.�:c�4�B�_�b*c��D����a�[�^���e{s�K��-��֦+f�U�_'I�����g_\�9�?�})a\+$�4����d�
W���_�SZRp%e�"�F��}�����Qɇ��9̖�ҍ"sbOz�R1�T;y�`�׹��{��P"�l������b�{����0�v��i��n�ܥ��;.�d��@�����?�.����]�¤G>,8�ճ0�M��k�^�Cbf��{��(��=$�}��fJi����Y��A�c�\G�p�ɼ��&��ʲ�e}�f��c�oj�!��M9�mRBԳ/�֦P!	����z�1���Џ�;%�/�\�ݟ���Y�!����K�m%
�����^ȷ+���:�O�8��$���N����Ԕ5��q�9^-��1�~\
�>�>]ǲ�j��2W���6��}�g-pP�<7�u�h` �qŽW���7������������X�7az+�A��0&)��%����Ч�u4u4In$ό4�g�ULhLT�*bsuppj��ڄw�¾�c#_P�,j��6���~y�0j�p�(+�������q�W�{��8 <�ۃŝC���]@kF��q��uQQ�JJ�H���1���@���Z=��֠JS7��ս��ZO�8R`��~��̣�ڃ���_k*�,hS7f�z�L�~<��/�<w���T"�j��8�NX����A(�Dd;�%��xx��YC�zi� zN�x�L^����	8f]1Πm���5�
˲�;�o.^�딻\ya�w�)�,���24rQ�7YKg[	����˽S����!�S'#Љ�=Xǜ;Y�,�0���o��vH�6��7�<���U��>C�,���M�KT%�5-l1s��dn]�����Lz��:�/S�&���L�tt܃�Ĥ]H�1�@\K�������\���W�"\<��:��6���a�W�d��ɾ$�V�X�~�hh�_6=�K�1��o�^&����N�F�d��XY�c�X�g|�?����Ԩ
�u�q�N	����U(%ޢ������/ ��il!b5|;N�8�1�_Ǔ��*�kҐ�����ò�MH�%� Ő�C��Ǽ�p��A#�����n���~�>7_G[,>5�D�柍)��h���ϒ�;@�f���Fs�c��xE����Ӵ�E�
�hxs.zy�ZF\�zA�'4�_��Ϣ���.�OԉN��uq0�"33����2��r�[uNj����ԏpГ���B�t��'Ϧy�*&ky##3.��G�C��Zj������?�~�a`Y��v����}���>�|	�H�W��I+mL��C��,ܫ�T2�'' �߅:y�53A*�a�j�gGL�$"]��������1aJ��U�'�W���||)b�_��J���"�\CR��~�x�������3�$$�Ie~�$2����^��Z=���河G�5��{Y�N�X%BP���f+���K!��ܘQ�@݋�x��V|0�>��R{[E�ӼZ����By3?���޼���2lKXإ��ߟ�;1Z�Y�A`��r�=�-M�m��ъB
Phk�Sd��1������>�3���@8��aTu�%����q#�4�>�m�
�6����)���s5��v�72CfC��<e����}9��ψ�Z�y���٢�J�V*)ڱ�5������;e"k��8v&@��*։�(*��ra4�_T�*�?c��A�|� 4�T�y����?�!���Iew�T��8K'���Do��[��4B��A:����6/f��'p�DW�^��kA��^�Ԃz�A���c���e��VU~�)��y��&(��C[z����� >η̂���0��3��7V=����)N�[;43~�z!��C|��A�u�!�J�,%�'��Y���\��p�P��F�m+��L���p�����Zt��0�����q�s*-@٦&>9�.�=R���w���ǩP�֣�?�ll|���YH�()��Q*RX�4�T��("�"n��^]�G��y�U����۱�~�0g�ɯl3����AY��he�~�6��#����g���e�wa4�~��m5�6U�q���=���я����O��,�
 n��ʦ�j��Qm����f��\��=K��x	rHD���[q񏋒|O��&\���ј	un�Tq@i)�B�c���aW�=�)��l���`��2����
z�S��?�A�$���{�6Sj^p�a�e��p9�y�Y�b ���i��y��u�m�8N����:֡�I�z;�*��/CB�,�l��� �Z���dk#3){c�'�}4��4j��!��d�+��l,������]�е[}(��-E�*֛��-����ˤF�*-���)���P��T���p����:��q�AX��<E#� �SkL(�(�j?}l�<v~�TRU0h\��+�u�o����(JlCMus~����r���]Z�J4���;a�ۤN��{X��S޹�ov��'�\B�r�*��|������]�)O$�1j �(�duY5ݩ���Ĳ�bv�;���R �� ���	�qv�0��{�ҹ��Ąt�k�$�<�32+�U24���)#m�fd��i��9��b1lO=�D��/>��*O4�[���'�l������r7�%�u0�7n%!<h4in�aՖ�s�,d�������
�맭��w��wŗ���5p=!P���"5
+E���tȗ]�Ar/�����\a.J������OQ����_�f�wmQ5p�1�)�1��P&��,��N�k��"2g�'܌;מ��>wΚ�� �#B��.�u�Ygݡ�8q����6{`;���qb%�Xa���
ֶo��68{=�t,p��H�k�)�$���D���ͼu����tcc\@�U�f6w��|�.�iFoȻm��@��4Gi1b1��T1�<u����e��E�������44�LwNj!�o�Vd���o}*-���nF��[T;�����}���:��*��W�H�1�F[�K��#�,RC��G�Q�M�vuN���N� N0�H4h�uE~�o-q���Q�C�Չ��<�p`���u��J.y� �=*N�åA�C�^/6�C����Vy;��DnJ{U.us7����I��w'H�ŗt~�٣x��aR��ydq�MJ�3E�A͗?aHV�||-�J�F�<l��1qt�l%�K��(�M+�l���i�P�="�dF2e�"ǡ�n6��K��&Z���-_��ʮ���e�D��-:�E_�ݾ|���?���g�h���i��wuJ�zS茼w6�>7&���44$����Yo��U�+�k%ڃ͜n9ʨAE���T=~�@�V]�S��d��S��$~p�^�^t>��������c��`��u��]ii3�P! �Xx��I�]�/�����I1���v��$�P�a�pi!�1���J�=�O���8�2�v��<VQ��-�u|$��K��
�p^��Gz�"|�c o�����d Dʠ[Q�'�ř�?JM ��V�G�\����D����EC�j-OcdC�]W����o�&�4�LO���(�D�9i�>���r|l�����bj����1�c�g���2�జ�׉�HgU?\��P�ѽc�����_�Ұ�
�b����0��ٔ�`���Q<Mx h��E�l���d2��u\}���_���(z�wp�t����	hܥ���N��%�s�&�J�����v��T����ap��cݫX��7)j�ܹ1��xl,56d��)~���=n��q	�QR��o���c�R>]�!ټe�9޲�Ƹ�S���h�i�%9�8�Dłt���xF��C۝�f�-��2�O6Rz�?���t���$��3�xMA������@�*r�	��0(���� �.B/��VO�2�-{�ͤh�h.��x�b
����+�C�vN�fM@V�R"���	����?�(���%��>1���5���$���ݦ��v��N]�