XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������C�S'���-Y�r=29��[�;Y��2}:#qK�+�����+$U6�C�c�9����z�΂���0�e�@/��L,��<k��I��Y����*��{�Mg1��	7�V�^�y{0���PMNIO(���Y���V/.1����d�dǑ�<ch��q���lp��f?ZO�ѡ��������\"��|;�`���4~��d�#r�l]���ZÆ���T�q�L���m�/�"3��O_��B�)s��~��f9��`�X	wK�C'jl��>rHV��v�-}A�<fQB�)7��7��a��N�#@��#+�����o��L#5�b�J��$���w.�3��AC
@��t�c�(Ъ�^
tr_��������Ng�:�W܇�P�������j�(ul���Js�z��e��>��*���S���b
[�ӗ����w!��K��-D!���!���}����4Q��瘉,��IE����1I9s�#�"~Tb|�ן����:x�\%�������Ej����V��`���U����^��#B�w�F�]|zМ�DE�:Ou�E���e.&N5�7�]�E��	��|D(+�+��B�$��r�����5�~������VC�m<�#�-��-�+��r�~�
c��l�l|n�JI�����*��|
�.-�u����&E�ȯ��$���r�$P���&Jn(�Fq���Ҷ̰������0s�y};|v%9���М!8��S���XlxVHYEB    5224    1740�i�ӹf����>������-�P�JХ�Y��<S�ri#�A�ծ�o������NF�����#�����@!�R�>���/�)z��]Uĝs�	�6D%��Td��-g:�Y���3���|�� ����F�&6���O�!��Km�j���^�������{���b���g��rb �U�~�W�[�Kb%	�{%7�k�N�;�	u5�t���@F8ݲIo�Hgs���� ��	?
z�w҂���{=_a{W̅5⨬bZv"?*�,wl9�]��x12���~���k�r��v���M�L��������$Y)��������`��s����0|����N�i���)��df���w���2��:RA'��K�L��@-�*T�X��F�NP'��;:o�&ۏ��>!i�C���t		6r0M)$+��sљZz�P��I�e�)��g��GCfƶ�Ϟ��2�ٹ~>^�R�;��������Z���a�Vk.B"�+t�g?�̛u�#��n���.j/b����E��a�,�Q�,�4i�e[7��;�F#���eG��@�L���,�� �b�J�K�����Eќ#�䥤����7/�Oi����	�[Ѱ�o��m�u�~��~n�P�[���d�l��`�x�wN5sKG	Vѣ�aM%,�px���>��i�1��}���P�k��z/xΧdo�6F.G�V����aU����2ͽ+�̬�AګEqINIq��f5�I�r](�^0N�x
��>N�]͂����8u������oJ��U�h{�<�0jm`淽ν�����$������� �v6�9���[��X�ƭ�5����a��w�	Ew ���̴,��EU��ʚ�9�Ю��J����^����[��PwU�u���O�:�Ճ9�����7pNNk��0]� �48[��9#ז�h�6L^�;�y���ѱ�Ĳ8?4�`?;�����bp_?�:�T��<]�3#�RXȺ����K�8D�+f���=u����^AN��\�5%��r��D��x��ҍ�T+|!D&�ᵜ�OHɶ�;I�I��윓�Qt�ir��&�8���G�P<����ߣ�;�-�f��sp������4����2U��OҙD��N�N��ߊ��5��V�y���#�Z���z7�������ཌ�:�a��L?µ��8�V��%��	�ب9�	E�������*Ȓ毴�t� ����T��n��j]�^�֪n�'�d����#JK��}罐
f.�η���t�w�Q�Sv�b��K�4�Sk���'t�3���<ٝ�������r��Q�|w�2�O�Oe�&(�j�WTY���(A�|���n����q�mpɓAW�όx)w��.�[�r�G��-t�"y���C�߀�p��l*���g��&�TԢo��E�ίÐ������݉{�V{���9��eѽA��Mz� ��'�7��=�܄D-��
ɨ{� �1�º���q2WsM��|d��&�ύ(ǀ#��3��<�����yXyY9�ϣ���,�ϭɏ�����
w�x-��&�v~y�
�t���Y��^��E�jp�ú}�B���cΉ�V|�Ws�vْ`���yS��n�x�x��1�_��91���;�*�&炢频xΝ�yw}�����f�ܞ����g������8��*��%��p��zw���Hk�re���_Rlp�G0AWEK(v:|b�ܵq����"If��̥d﹙�׃����N60�]WV}V�>�8ӍH���]�;��}y5���'�;Q��7;�]�x̰�"�r��3�}���d��%��X���b��p��&���,,�cBy,����f�Q����/�[�)�������[���-��I� �|�f/������px:���5��4�B!N���Ov{n�{?�aҦ�:�!����`��k/ |�";-���� a����Y ���#�ξp�1V�����-��M���
f�W��i�GY �K ��EUh��ok���	�#k�����;�an���N��&s��`��]�Kl{8���)Z�/Rm����e87�F��
GPo�5�W�h�YP���G�Ř.V-8}�BW6��Pz���<dΫ�@��fVn�h_����`��NVĎ�TĪ% ���Ί��p�[�(��X0)��[H��TnI.����G��1�P�K�KD�ߧ��3q����%1)���|��Hڈ�Xu�/j\�-�u��o��td�	NU�V�
&�ou�-
�����G�*/7Xe|%,������x(�N]��!��Pd�^6ŒJ�#�������+(e�`J���ج����(]}�|T��KV�ޤ�nL�mC� h"+r��5Pu=*ԄԘ:�����8r�	����\�+I�\����0��rA̽^���;*\�@=Zi��a�&�����tR�k���SƩ�j����d�J	�SGX"K�5�'��Z}�ΫQeP�U����ܯ������l�dI�)_�v��q7vZwߞV�+=Z��C{-��,Iu2t�'�I��3��,�qY���D�������j�����@p��6����("K�� ����S܎��D~�D��Vό[U�ؗ���@��5Re���Qc���O��e��>�_�ǔG�[[z/$��<$>�q����RɃP+5ʠ�f��ᾔa��QH���"w�� ��hEBpf�&�ׄ4�%�!I
)߭���@Ob��j�s��Oc��ٕ��U�31�A̶s3�/��J�����ܐ��2��Fjs�6�p���#\oѡW&H�������>�A��쟇�e�?*�7��UYcG��a����V��MV��Yr�&�!�K��$co4���<ȯ1�)P�:;Ē}#�
Ge�@:$��0K��L��V���w�E��n�a�"@�.�L���#�TKЕ̩G�XN�I�QN�K`��u��Z ����R�sB#	o�	ED�+/L���`�C�����eu�AW��>����.�����r�M��5hg�6����o�A��8�w��.dP�s!AtP���J�3De�A|�\}�I~Z���&��@pT�zMԎ<�l����u�ܡ.ٳQ�%����J��ԓ���ڶ�P/�'(%E;�Y6�!/
��oY���<?ٶ{iB�}�*���@/(�ݏI7/��"H}"� �\
,���1%�)��#�T�g�����F��6�}�1�����l*�^����ΎĽujxi�W\?�g�M^�����?8u��YtN?~8�> �
:�D�KW�A���� �3Jt���((����}j~���	���k��I�����5�蔘�(�;#�������6��� ɠ2�]�Zt�E�5�Z_��3��=��[��)��ˈ=��^��e���T�h�Jku��p������|�R����^y�h!c��i���g��S��o�w�<�tI7��5�!D�c|��k;�����p� �����颺eX�i!( }�]wCE퓶VU1)]�N\R�	�mw��Y���N�2�l����8�gĴ�0ޝ�t��@�I:�����qm4��y���y,+ڻ����L�:| tá�\9��O�Ӝ�.��H�����o,@�A�0���Z L�^��qd�%l��TJ��u��Ю����vJx)�_���&�S�͔�ч锨�2���OH�2'_W�r�b�q�Ϫ��d�C�)B�K��?�x~oٻ<����+W9x���Ћh^���4�տ�����)Q	����H��S�,����e}D&���T�g�FI-�XM8R�E�TP�ӱ,��z�g��<f���Iu���|t�ƌ+V�R�@��D?����:&B������O��z���ʢx�~L�?���)C���ju�o0P���{�	��� �����$�wT� .x3��i��)�3ү����)�-��,>8���x��M,۳��M?�G�NT#�W�֍R�˪\�d�9��0���Q �PU��+s�ܛ�Dh��8�)W|a\p��8�Ob��~�x[Fl�Ga�E�#d�9��&�*�S,oP��A��z�A�2���21hO�!Эj�bJ��B|�Y9M��	��/���K�q$5a�H�7UX�����h8*W��AL4��u��kS����X���ZH���-侳� �V�O#�"Zm�A�C�7t��������n�Hb��׽Eb��O��5����_e�`)D��+�ւ��6�Iƽ����f��T
�$Ʉ�N&ŊO�n�0w�@(��{�őhˉG� ���<Vv[U`�� �w!�G׽4�-����%̜�e���b�R��T10]}-����'ڀQ_a�/9�#��Wc�|�Ԗw�%�/��p	؟���*`��{-��(Ɓ��l���;���^��}���u��Y����p�t'��zV�2h���ZyvZ�: ���"�Gh��L|oE��)E�b�᳢����B@��1��>E3үTW��\��ﻕS|���A����Sl��=�dW��cQ��̳�B���1�#������]-]ο�ye�%֒���]�b'�{c ����(��ʧ>?�<33�`� �(��o�@H^�F���_�h,̀5��
���i1�xz�%�^�,W��Y�5��&G�R��[�������"���s<t2�)�8-� �����?E���<�fB��ஜ	�M��Pn��6�ZBI�����H�H���Ɛt�j,��o�`��2b(V��o��
���x3�P53���j0S�#��2����`�Z�[x��R��+[�~�Se]H���ck�8M���'�X�жH����A�cI��*��t�mr�[z%�0�E�#;��ܠ���U�b��y �N�������ې0)}E¡�+�TpKYO��pó�x%�Adnn��M�Tw�������チ��r�r���q.0�	ذ�'�w�o@��Q5�>c v��D�^"P)g6��g�l�t�� ����w�hE���Ȇ��S������y�Kɜ�����&��M�,���>E0YO��5ȳ�+E��vsd8v.#;Rː�V�Ŋ|X�����aX����q�L�<[�ㄛ���XjdT���7̷{��-^h*�E��7�}�p?���P ��{]�yׁWēD���C���|�E�g��(.�vV�K��`�����N�=�m\���q$&���Y9Y$Dľ�%w�ߐ���B�XM ��3evGZ)�z���t�������F0~���B�c'K9�PC��{YlNo{�L���.'��ƙN1��y�/�Ҁ��?Jy��A����B~�i�z��.�x�����@q����ul�F�@}9��6��SY%�!q�8;��`N�\���`;7F[e��Y���6o(�~� ������)4�5m?!&�(C0�܅��a������z���n�l���V��<,C�o��Z)��d��~6DV�4��� s��yp|�1&]�e��d�`'�f����POd�sA�/�d����2Ԭ赃R��J�A.]2^@���<n�r3��@>�In�}hP)���*�(�p׼� �����ӖS��غ#�YN�þ���^��.j1)��`�uA�wFgҖ���ҡD�^βݳ29��� X0O�I��U�5p�kQ�5׷ZYM���/�1�$O��יKtT�0I�?y�An��l�pq�2��Φ3���B?�܍sY]�d%��ۯ82-���ɼ�װw:F����~J�l�������O��`��L�; ��r`�	WoCfQ�=
R�PU�Y�)�'�~	i/��� ��Q�K	ӎ�U���U>�+=W�j�D
��k9��Ӵg�:����o0