XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������n7��<J��<���Gf��gҥ�;Q��hÑ��LZ� =Ƨw\��R;��P�Q�r�� ����
�ڼ�<��_r�a�Fq�̩�
3�A#��F=2p�Z>�`p>$3����(i唑G�����\�+*����������o9<V���O-�e�0���8K+D��(lE�ټ��&,$�)@�?k�>�^dS��p�r>�:C�UC��#�f �C��HQY��q%K�t�����P^u�'��y|p�uhO9d�kA:�<�6��O4|=�%�����A�i��=G'3M'������xݭJ�Ę�Oz��$�c���E�t-Q���:Ͼ	\Si�&T4�9|Q�{�n#\�#T��pb���%qâ���n;�c��s�ǀT9Iy���v���'7�����F��Gg�RbWYօ H�����������j����Y��T���"Pz�n�� H鲁ᜳF�@!�M�b����k��%��.�"�!v����Tq��<DQ��D�m�!k�k���O�F��J��E�i䇴Iu�8�W`$�)��}ϧٹ�&CA���-�a �	Ʀ?�bf�,�+&k)�I�*�y�A���и_>�d��C�]ܵ�u�{=�y���Y6��iz@�<���v:wH��4
D�h�
�����gq���v3�	�ި0��Un��_ cP�
noU�������A���.8i��*�X�^ ��Ku1�T�|sD��VoO�S�V)�y�z�?D��Ev�@��o�3�XlxVHYEB    39de    1170JU93j�����2�GtZ�p�A�;�/��ۑ���v���>��MJP�h���H�V	�g�m`y,��ɢ��:}������J��Z���2��M�Ք�m>�..��<��|��@b�POGp�L�7mۺ����
�3(��>١?�-������1i��R�8�o��%�%�[��9����p�f�|��P}�,�v(�F�K���o��A�ߦ�.ubh��q�bQ�W�����ww���$�MTsw�2� ��xs�`���^j!)B^q�1JV(��E�!���n�T��v�=B��������Բ�l,���}�O.��*Emu����w0}돥��W��ȑq��W~��h#G����Q�����ջ��R<�v+�����Sv(�ؘ'�'��u�F�}����� gb`jhs5�;��Q�H߄2m�1�`Y�#F����ob��>���ب�F��)��	����*9u�L��X���3Bʈ���G�i���G���{K|�����[Qc���;u���"�Ҹ;�|�|�Q*�{є"R�7_����m�� �SN�_�c��{b����n�<@���z��IJ2{^g�</p��zy�$�7eȲ
W�m���8�f��2Ҟ�
�;8{��p%K�nqN��G�f�[k1�vua������ҏ��4eE+�:��uI��� Ni�&�s���D��?d5	h���-���o��L��|�@x�
f>���@Y[8�n�9g��{�*B�ma�C���Gb�P���ۏ���졿3��sd�.e&�)���{u�!���;��Ί��'�Ȭ0�������~uþ'����b{�#����w�'��w/o6��%u�Np
tE	�kʂ!��C�J#Z�A7�MG~��H'�t���hlx]7o$�X�������m&���1���+���S((mG�C��&�}�����ăP�a����ξ��R��@Y��n�|ٲ��,ٕtPg�,����w���AE�(�d�f���z^b�O�E�&U��ꄢm0�>��"�L@8[�
�nqӴxy6�l�$#�NCD���&R������Jz�b�.ђF�[΢.G���t�G�a�eR���L=#�;��l�R?<i��Nc)��Μ�bE�W9�;��ޅ��{��W[z:�.�>�h9�p@��X ���wTm�F��`�T�J���K�օIH�]�Ƞ���	g]�����-	~�ŧd��W�F��D���P��x;+p��¿`�N��7�|�K1s|���ÿZo^���1�A�����>�~�L�d��Lop�-�廱�+����q�G=��_�nv'ؘpJR����h��3`��wĦ	d�kt0;pŦ���I�G���$Pj�u��E`�k�q[�V Cۭ�\�K�yۃ��^�q��m�� ��|?-�eR�P�5'v4�˓�Cp��*��@�k|��|w0��J�b|���mm��.*\i�k��N#�'��I.�oz���H�F��t�%��i�T����	ũ��A�@u9A��+��1=�LC�j/�Us�+����e#BWnL�	��T-œ_�����7�i���!��eS>q��g_�"�`ߔ\�Q�X�r|�թ���4X�#D`����p�g������ �[V��ʒA�UԿ�`�H�J���B�^�i��@����\03Uz���w!B�� ���Aw
$�4G�|�����W�������!��1��5~;��cz��|剌�yO�i�����&��p%2;m+iM�92�<����ϭ��.��g7�����7���-w�s�L!�7C��3�K�o���I�Y/��v�e�C�t�/ǵB�� ]\��$*R�K�V�%���������#�2Y���P��f=�L�?���z:���b��`Gg�#p.0��T���B?��/�������L�ͬG��f�sS�� �"ǥ���3c�*»W
���yP������v�=�q��{�|N[y�K�V�뗌�_=���5�M����p|߱�[kV�&��p7�]HHT�<�'>����Yd�M*�[�~)\���2����;�=��W�i���3 ��Ѭەi�{|r��s1��O�d�՞���pC�4���!����hG��h\ʏn�eRN�O�Y��?�12C`n��(�E���k�ß��]�~����@C~�Y)���� ��y]��W��u@��~{B��z~�>��p
�(�T��ja��Y�Q�Q폃GY�ʿ�����zݦg:2�w��?���?=�����`�$PoZ��,B'����nGB�u�p�{Y¾ �:�o��a$�P�4*��mH"�e��!/���0��/@��V���4�D�lW�jMr���i��#O2�`���[%i4�Yɿ�ŕ<(��.���(t=(��U��,w�����e-��%�m�T���W9�)�,���e�׎=n�����$H�C�tn4$����[.��tMɺ��t� 뻏~f2�)�e��4-'u#���me5���6-�_��9�`��g��Տ��p+����_��j�poYP��;T�pf�R���.�;%v��ZM�0?ry�c��O�K�o�B@�G��� ks1�e�3�t�c�w6�焧��i�Ttin����G��^n��f|���+�b1=���/Z� �����EᏬ�%�}#���N��!(+4u���Vq�Dޏ��i�70`���IO4o���G�P�-�#�;L��)� ����z�J��  �u�K������=���m}����E!ܵ�?9<���?p�UT� ������5,�I���4�+w�� ����;�\=���G�9�g�!؀Fa<�ʾ;�)���|�Y^q�`����.ʝ���5�Z^�\�c��$+��������`�5Y7`�/��R����F��ZT4��)��}.Ma*�K"��A<��&�� c3�黨�VTXp{���Gm��@P&�&8�#MVM.�wz��O3��N�6��&{�S���=�9�xx�]ȓoB��E��^���X�.	& ����CQ���Mz��bV��$w��iR�%E���}��nXO�q��i^��f���Y�`n��:w�N,�]��cα���_�OY�|P|��(�>ӣbxs�x|4��c~��']���oJ�G�E�-{��'a�(!e���R���+k��#�A�zq��UPԺ��Wvw��:Al%q1� Q�0˕����0o����װۘ��,���{B�.���(\���}5����Mf��wD)����-(0"
�?�l)������<�xA���R�]��~�:�������rfG�N�I��ZF�}�����K*`��<��q�C�:-)[>�>1���nh��J�@����0�ΠBB2�Ȧ	9VT�r⛾���bR�ᡵ;e�W���h�d)���%�R4Վ(3�d��s���;��Մ�����4l�~�V��#�ʉ��$��n��U�W��ok�¦pi���Ѓ����y�ӽ��а�w�D�&��3����c�΂Y��g<1�x�'�{�E�y��7Nq[��^dO��]GTȺ`Z��\��֚��`:��x=����H(��eQ�	��.�_S��k����0@����t��I�䓽�ܟ�nPh�ytN4��N�jWx��bI�F@HZ��gFK9��?uRQ��gI+����=� ǄԜ�K).
�%#��h[���-��<��'@ܡ�02xOq��ݗ��/�[?t�����J��x�R�a�,�] �,	&�����������[z�x�3�,���`��jR� ԯ��:��l�@x^����og!ۏҨe)�$���?d�N9�"� �*ॺ��IR�+Jv��z�?�f%5�&(P���u a�C��K��]�h~$j������op\�sC��s/%L��	�":��,�[q(�H��Ձ�	�@�l�8���,*lWy8�c7�u��ђdu����g��c�dXaʌ(�K���@x�7I��/��-�g>�]��굀��[K��%�%��O���`C�� m�����{�Ajkg��ꌅr�t+Ŧ�cO�96%�SHG�[������1$J1��	�� ��8��I����\�uGx�d��%j��"��.(���f$Ჷ�]�ߙ�R. ;���z�@�W�A�Y������2*�8L�z̀V� P�c��_!D�y�+�����|��i-,n�p��$�:'%���:,�=�34�{sP|q����T�f�ң:F��z�m����F-�-����Թ��2��� n����%v'����_�H���w=�Sq��iu���U�'XD|�q6_]j��FH=^��)�R�#fЬ4�;A�7�l�W���-��A�ըa��z� 7���\����³9�:�������c