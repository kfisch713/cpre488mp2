XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#w��FU�|���R����8˷�4��dТ���1��7�7.�K�v����ĹZL]�-���&��P��O�[��b�j�.}�V��"5�mꡥ�y�sFé �.9���`�R<y���Pi�υ6y�%xg� ��.+F$�_��]��T�U�~��(�}coF��Er���E7�&�8Xk�b-����	��*�n^����{\M�̳���x��$�-��M�������3���*e�\�Pȏf� Iw5��c��>�Ga�D;!*ؕ��OH6eΚ�w��%�+��=��U��"��8�������n�N��0�@Z�\��&��Y�1�PIz:|��@���:&���EdV�Rh7?+xT-��v����\����?[.: ����g��l`�/��.5Y�]�y��B�]��a[*�(�a�0�h�"��;Y�}�1��)p���5w37��Mt*v���W
�>�%���D�0�Z�z�Ki	DZ�����Ƶ����P|h��eEB�����Z�8�kɣ	���1�ha��o?��L2C�Q�d�*��-Un�\[���a��|PSo�Js�6��_�I\�/AMl�p?C��*0&��,�b�C1�<q"TSD��g׻!��[l�v%�{����>��|���H��{���^�=���.O���x|&�C|�Gh0x�I8H\�[��A��n^~�����f�
(0�Ff:�Y�C9�A�A&� s�@��N��%�C����T5��GFH0Q��S�;iXlxVHYEB    28ae     b60QgrBΞ-f��#���֍�� ]��T�,c廋��w�ZWù��������}���D��w%�m�dc��lP�х�ٌ���ǃ���k$��2�~�_N�ݭ!14ϫH>�x���5*ţo��?��4.�h]�|��E��
��&ms`����~z��W2�k��rd%?��� ����_׷���ǲ�n
��h8q�w�ꕯ�ʷ�����}v���
��P�Id;p��85�ѿ���Q�h��Ő�nM�bfΆ�^������Y�����G�b���Pm��ږ��g�͌�H���<@��h��K�@,�2���ݙY`}X�t�0V{ �k��>[uy�K�;%�~��웚�0����e;
_�PZHFv�JE����t�d4�];[�j��AFx��+�ɝ�$�w�S,��'�� U��̩�q�JS}��G���dR�iQs�č`�j�5�7��#��,�-J��V�A��g$�_�Ѧ5b{��#��׎~A#��wĥ���̍j����I�X�M��yG;�����]�P��~�T��f�hu@���ʑ�p@w|JxvKOLC{�,�ҙ;6T«�1r�sN@����A��*��TK[h���ݬ\=��ג��(��b��{@�Hx��bڲ\�Ak��M�H���� �DN��-6~y�77w3�.��y��~��t�Ď���~!��/�Ԣl�~�?[�q�MU�cV���Ԉ���~Q<Lf��'��'�
�
�*���38�Q�_�D^ ���R�y��WA�FN��l���� PX���ߜ���{1q��i:�͚��W��),b�59j��|$�.��\�֋a��"�T&�xճ��s�O���|���:y�M� B��E�/ɂ����V�z#�3�E���;4������������{eI�q\0x�]Jt�bD?ˌG$bks� ���5ӛ͘]� e��� &�z��I4�r�����(��-�Na{&TO��T3b��e% ����h/ٶͼ~|?-�7�?�o1eC_�����Nu�n<ӝ
^��=I���[V�="o����@*�����s���oQU�Xͣ�E��{)�?m���g�i�A!�	:�3~<bwh־�ɏo`OZ.���"�؃Ry�ȏE-^���2!�n�=#��n�=P�Of
Y1,�"�k]�k�a�Di�0�����p7��ͯ Z�hR_�k��P�L�a��#4Pb�
��iċ�gO��7��9�θ�8���J}0n���5:FI3�ځ��o��lO��Ȁ�L�:Zm��$�TV��C�l+���*�sq�me4�V�U83N����ɨ�$my�/�C���J����tF5D	�P�]2�T��o�#��l��Y�u)�1Dy8����O�_����W'lՓ�8���g/��j���*���׾e�)�sǩ�+�)�V}��| �-�~�|>�k��5m�Gb��(��� ����h��r�#)>�����P.kǘ^EQ(�5�XK�R�xzp$h��l�o�.`�QxO��<?^��3/�n��q�:\���a���T�|�`!"�����
=�π�
h��"�t`zd�%�QP�Z���t75�e+����0�]=���Ff(|�������q�NX��$����8oCd-ɱϴ�L{y��+����`��֕H���|�Z$D#B��J�ҬCK�ha�ڭ@�a����J(㔶|��ܻ����7�)��9ƙ��}�C�	ҵ˵���JT\�F���wv��x�|a腡���>J[��~:	yBO���7��+�c��=�Y���O���p��ǜ��Z/�/(N�i��#"�,�Z�F�mr�_��
[ZN���b��O �^ 9�1��	 ��+4�y�e=s	ܾ�#.���U�OX�[!��O�m�Eg4U�,_�Ə�����H����E������b
9����^�wz���V��-���g���y�$*MԅTq�Yp�행�o�j�������#�*8�ngj�����'�stE��V6� 71_�������2���EU���c�^yq��$J�hq��X��O^L�|��9k��K�����B9�
F�n��0��_��HjG(1v�R�cݣ�ADq�j�ͦ�Rw�'\�;��_e��7Pn�S��6+�5��.����Ef���Z�61�WG\��t�s�CM��g��#ܵ�a��ƫ�$����qwN�>n�}�.�
}��r�-)�<F�=4�v+�}�]{�I����q�e��!�$y�ʴF�J@9+~�o���U�:��턽8����O��iV���l��t;��+��N	p�C?���~��G���7J�c�y�Z �G�W"pp��y�3�������(izaWCf���}�+p�5���a�/髷��2��4;��O:�?܍�6��V��d�_=�	N@�	F焊���(�c�8��@}�#�A&,Z媽�R��z=�i�j����(2�b��Zj�~��5&��J2B��>��=��k�����&㎄�_��U��(_����v�D���6i�<��y��#�c���~��֋���w=��5��dvA6�fP܈
+��q�S�Nң��L�����	�0����˼�*�!v�Ys�4��~yh�TT�9�����GgC�QqT��f%4~ܶM}8���=c����#���$|� }�x��27�q��P��Vgi��Vs�kb�@���m�������)�-���b�`c4,e"[;�/�<����$0�Y��aH��¿�]k�m�Џ�)*ްW;m��}J,��3�,����ڋC,8�'l�$��.�^k�FdW�7����,����Ռ�5g���p3r jֶ�`��~-;Q�յ:2|�n�%�7�