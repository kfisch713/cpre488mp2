XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I��Q�*	A���;�Q��hx�o����%��h����c��a��A��Afz�F;\��/,_#@� 0`y���%��|\��f��ȅP��i��(���
���r�_εu���p��Ϗ.ZcZ�6=��͒���Z����w:��i����os��
݉��K0�qH�4�O���pFk��Af�L�5;���Y(�(E!��i���}{eZ�8���8/��#ܰ�}�Q#n���2���Ң��)j�L	=��8�����j��
s3VV�7FȽuh�x@$��fEHb�c�o�`�jH�:^�ۍ�	�]��|����.�z�Ln�m���]��=��ah�bcP}�.���MzT�o��ȍ R`��ӕ��hk:D�N��֫&�@f��wXD�s�,���E^���Y��d4ҕ٦�Ӻ���Y@I���k�;��Z�d�8�z�I
~/8	3��_�/��5��F�tg�u��a����O�r~y�� �
�!syd8��m��O;P�;�;$�+�B��)��FN�Vd@�P	,2:a���]����0!��Ýl 9х��D��\r���l}��ŔҾ^���O��ͶJ��׎W�8����)�����2(XD��S��]}��z�O��ƻl�6�n�o4Rǹ���G`;G��}�~w�]xp\wr\jƈp�셺q���]"<����!����Q�y�܇�����7$����!<�&-����&�k[����{Q��tR�;�7���~��wXlxVHYEB    dd8f    2160s�k{ S������˴3oi�L���<9�}��3���k�*��l&�v_�Ԗ�Q��>�Y�����U����v�|+,���^`��F�]]͡��'챺J7�U��	qzV�>�m�u�z���b9n�é3xU��P�gi������#���K�7���~���ۀƼ����1�Tu
�W����H�ɱ�Z���6%��r��*�@�Wyޘ���x��Sۄt2�/|{GK�M#���ʊ�=眜h�>����-������\X�^ڜ<G��nm�XK�Z��Һ����[^��g���*�\��o]&�,#�S���x�&.��m�>�G�]�H�d��5��4��<(���d�k,}�����@����̚[�0]�Z�G��|`�s�����ԮKJ}=��Q�93�p�|g�I>��.ؖ�z3~���(/�=�h�+�����cLr����{�E<0(�9��cX�&* �=i�z`�aYP�
L��O'Ҫ�ཱྀ��C�a�5]�����l�ɽ@���r��x,|J^���nо�D�t�-�)L/��x���4HR�N,j�n�f��;w�+,�*|�DW���^�S���4oV9�Ǝ�8�䜫��f8�h_��o�7:�e�bu&�p�2[��:ņyk����0P$1g7q-��ЍH� ���L[
Ҽ���XA(e�=D�[S�P�Y�2�O4D��zci!�"C"��E�B���)2�k� ��É�N�j�#��h�k��׊NfqN/z���#�G�|t�[3�L��Z����X;���պ� EU�&3����as��~U<�?�i�Ӡi[��=O�ǮLh��٣&�i��xBj��S�q��qS���ff�X����"D��@hx����/*�oD-'��~����*,���K�6����1�	���Dd4�+S^���������\p8�2���_�c�<�`��O_ X`���[����t�fG(Bt�bS�L|�s��	|&�v�w>�"�n���[Ҍ���Is�ۜN�Hd�!q�����M�������?ye���y��C�p�<@����s>R=@�|��\8��1jp�Ȥ�:{�'?��D9 L�YUYk?�sV5��DzFq�-WgQ������h��ri5���݃{��N\͟5���Vi��϶�L�־�&�[K�|��QFI�F���������{���4�;㆒r�{P��>�%���I��{sW��,��o��K�z�Ი{*��n��}]�:%�R�X]�')	�"U�l��M���]��=^#ꅘ���I*}�죂�wQ� �<}E����ʬ��UHW�K,*pn�������������o�V�j�/�֐\�c���.5����8�(�� ���xU�u}��X~�V��#����fd�vi�W��mYNǕ���~�\��q�r�HHy!D#/R���p���s��2=�rY� �J����h�9�I٤�q췅K�?A�11#)���͙�;�@h�B�N˺;� ��"A��C�
�\`[�n7k�\���"�:������`�p��w_T��n�'LL	A�����ǊX�h7�-�ȝgԥ�F�v��aU��Vu��#�u�Q�B�WB���x��e�w���4/%����NGv�����P���J�ن
����iF�\D_���m�N��C"�&k�
��Jzz*C��ѿ<���ə��HD����FdΕD�&��q�SXNǕV�-�j&�ә,1���nJ�����������ַ�k�J  }�8�W�JD�i���ϛ���N7��l/�J����z�hg�U��p��67;��7��T�A���q�8��������2� L���Z=`^2�P,�\��N�ʧ�6�9�U�Ⱦ)�� %�*B}	�K��.F5%��*'kD�zf	�r7G)nMp�.`�+v��졃��g�i-�J�<䋽�|�W�B�=�W�Wri���I�e+"�UR���ރ�x��)�\�x�����.��k)ѓ�L2�����'R"�Q���+�ϴ�^�v(k#��|���w�|�{o���� f5DKl9��ɿ�֩=��L�4NT�#Ց����,3�]�q~٫��������w���Y���.H����?������؈:�zL��H3��w�4xE#b�է��͸�{�����aۙ�X���@�<���I�_W��L�{��9���.�>G��<��T39t���i�Ϡ!6eEw�>,�s�!EN����GO�
ʓ�^��4N9̶������vy�=�A}���0���6y�7�?<E]f�=*7�GޜF<�eڗ�����N�3ܱ(͐yH�H��Q�,S��(�����J5���A8w��iV8i%�_��v���X�E�3We�\&�R�����Y�/����BÄ��c�jz��u����tM��D1����:E||%!���X�@g-�Y�my�C�*tOu�@�}LN�^��o�]>��Z?�6�N��Pa.�`�R�Ai3V��c��MPC�$Y]wC�.F��n܁���g���K|��xI��2��6g+���r<^G*�)4,%�H~�����I?�]�8��_{�^��
8��z��o��E=�� �,uս
	%�M��G��L+��.�6�A���/�*����5��iX���;�ek�,?N��9""��o�HGj�G����Q����-K���A(k:��bČ�g"d�P'�v��S#�n����v�C3�d�ܨY�����;�^�Xx���irp�=���St!�]�R�g6���@�j�LK�ܛo�w��\=��Z5�z�N�D���P�wd�y�p̭Q�#~���pֶ���m0��-V���j��]5��4��uɹh��6z�J������FJ�S|���>�8lbH">e
0G[S��&[�!��td��u��0e�)��:Ζ�#$�Nd�A���Q���!�>&�ˠ���M���4����u_0C��L���9�����dk�f{����Չ���C �L���d$ȹ���Q�6L�@��r�1&n�7��.s_���㦉�8���$m�X��P��@�Eδ�P���Km�WIZ}�3F��4��� A�vi
�o�)�T�U!���pƎ�zF��SQ�%�0�3��
���m�v�.��o�ԅ>%Zg ��3��Y �I�����u�j���� �������U���}N�Lȵ�⻋Xfo>b�n��Ϣ���9=N6��X@ߤ0*>�A�nŸ�nW�ߣu����5�yo<k�]t�����1�69w.�C/��α��\]w�A�����RC���C���Qԭ��V�Y4�B�g�=�z=��h4mI�� jo�T�!��t|�zt�b*f��V�el�U2�M,��>N[3	����	����?�? ��%T�*����^��CY�9���u�b(G%���e�pG�U�� ������/#�]m\����$3�N�Jd�����9Zcw�M��J�Ր����� 5��E�ߑ����H�/v�����ѯ���k�1687)�c��J ��V�H�zݗ��R}�"i��U�Xo+?2�49Ȅ(����1���*J�=�|��1��C``�0��$e|�
,��ޫ;Fe���h0�e���R�[�/۔� �v� =�o����
%�k����GZǕ��){������` �\�{3��i=�����K;���W��Bk�f����1��ppl7�ΝG�ЎEI�X]{�{��f�0X�,��]OS���(�pV-sp�k�M�Q?EH�}��O@��:{X�������zR����C��x���Ʀ�� ���2:�so��gjcJ����`wP箥GR&�X��2�;�q/7���;��^|{�h����S-��	q�>�*_��Mi0��v�J�Mj��
��!i<E.U)�^lG��!���$$	2H)�ѧ�K>�Х$BjB��D��ad�����<&��p���g�N","�(��R�!����c����F�]��i̺��%m6���_[��ۍ�wǀ�T5h���nw�C)�,@`��=����g�=^�v��Tʣ�ї�l~��_C��׆�����(�``����ݻŴ᱘h���ka<r!��TC���u9Ĩh�,<�;ھ���;~�oQ�9�v��D,N�K�_��ە��`#�Ϸ���јόĢ�z<c=�J!�����P-Gْr� �%�G�>7�����"`+%�
P��m�A��*�R�]�h�$Y���� �-.�S�-�W��0��}Y;�L���~PO������j-�y�J�OE�L��d� %�O	����1-����5+2PE����긪��W2��	˫��G��ϡ������>��ǚD]�IZ)�����������Zf����)�����FKU�J�@��x¶��,^i�x��ʶ�M�C�D>k��͐��X��d�wҧ�q(.��E���Z�?�"L��1r�~�L�@����rY� (�(_/��^W4��9�c���+aIq��e 1ڒy+!���M ^��NQ�Vf��.�Q�'�.�s����
�A�ɶ��2{�y���^�c���"�Z�j=ا��fސ~Z��ڠ��W�-�����Fc,yL�u,��ABL�WcS�L��GaU���0�D�$w���{߂�(@���V�;�M�vG�T<Ѝ6���A���� �g6�c�!Z����q}S$���J���������F����m[G��:�;@uOM��y�,���B�#a.�
����`>�A���P���>��{���O�Ѥ�fqK�zm�&ߛ������>
�@�	 Oo�T2@��\��~ ����;%2Η�[���,!���,T}���g����Щ$����'#�73~I4��%��zy���!ųX5lsdY^{��5_9<V�b����aw
�:=�Yf��(��)e�]+R�v��!�JJI���w����N�Y�.Q��)B��z��u��[ ��gܫ^I�06�]��"�]/.��Y�)���(�%8i��"����Z�_eӰL#GR(F�^CV�Պ��>Z?,������u��p<���%ɖz.�5Q���[�.���̾~n�x��&.9Ɛ�1^�-kq�:��rM��s:ٔ�A���\���s+
�\"�	��f)���ߓN���>d�'���OQ��F��Wt��m�sm�!mqކ��=��x�c���N+���y�=�"������P����_��V��<A����'�ఴUsf�(w��aC������k	��~/j|���No�Zg�!�z�r��o0�K���6�a��w��~|0�R��\��!�yί��������4h/���\�7�W�#OV�����8�(-8�&���D�(���'#]���Ґ�\y��Ln��-w�q=c̖sT�y��`i{6��h���1՞
��U�R� (���c-5MI�,��0��A$���j[9��f�
�-D�N�%=�+��Q�/���jb��a�����	���,d���q�ɼ�[#��"Fc�tA��/�~�����U�*d}0ǆ����M�,�e��Lؠٗƃ
�E%K���O���#A��=L���M��s�X-*H��I6ֽ�o���-:��|�=(�S�u�Y�����%�w�vL��Y����� �'�w<[�CoAؼ�/�k�R�~�M����.�~s.��!ru.T���
?�S���OH�1f��x�1�0�_��~��ȾGjE��()KK�RE�(��j@��>4�/��fa
��|Ъ����4�ll�2��P��w<���h�k���TJ��WA���RJ��gN���L�m�+6��t��$�QH[���+�Kw!��k{\+�3��ٹ",�`��%�ܼj6�wל*2	��C���y	 �zJ(�-Sm}N��܌F���ES&p�b�v��4��|h��_=)�4��\�u���: �x9�Oܠ�����ڥb�B��"H7�i����pqK��Y#�I Qj#�j�ช�5Y6�^�l½�u�'��ap�	QϽ�UHʸ�5K�]=�!�ťaMx�Р;T3�O�<Y-g� �?k�}�=�`����K� 6��:���k�yK�w��Ӕ_:i��x�R���շ�2ğM�*���VW�ƣ�ңe-z���o���$'/YÜN5��ë�=�/%��XFc�8���t~�w3f(;k�8)]I�jYp��s��Ι-%�!,���e":�
����vB�46�.7u%"��}�g��d�r���q�4��p�Ȁ9TZ�g�L	�ʪ𕴖j%�_b��1m0B0l��g��=7�(7`�U�������KP���o�F��'̹b︇o�yƋMR�l���P�E р�nĥi�O�A;�V�x����}%}���$f��0�������2s���\=�B]�1�O��6��f��Y�iмqA�T�.{�[R��z�d��`�`0ejIq���l}(�q-F��is37b��f ��qp���PHzL�'�$��<��ɪ����Z��Cv��9`���U�w���;cs2���y[�]/�����~�m�Cc@p�V�����ɠaA��vR�Y�<)�6�Pj���͈Ms�B���&����@���:�z&���} �B$  �O��{;�1S��i+|˷��D�*:s��:ՙg�L�#�,��b��[����{�OcL����\�]~��:��a��i�ɳ��E���	����1�����ǧAo J0�)"z�����������p�KV
#֪/^R�^���6��\V�C������N�8	�T��˗m��O�a�ץ����U#�Ү-5޴�M%�.��μ�(��y��ۘ=�h�L �4���Q=F�x6����I,�J##�?&�ѿ�
\㳷�
�\L��:�}�zK���~���Q:���xUyɨ`6����q�o�Q���^@[��V��?�&e�?'�����n����t�Mb�?���!^�e��:{	F�Y��Y��_���Y��Ɛ�}'g _�AIY� �.R��y�c�ޑ\J�� N7���Q Z�0��1T��k��0�4��W<�e��9�Pk��q��'�M�����۞�*H���}���T�z��ށ1>U���P�m�?��9�'��{$���G9��D�\���D3�Q)��)�#��O�:���'N7sW������;�~X��㈚�P�j
32QPS�`⽂K-��2�+�n���G>��@�Q��U�)G��)�gc��Z��Z���Zbhޥp��N!�9<�k�ES�A�V"�%:&�=t�rs�V7z�����w�?�?�_3F5Н�M�t)��a�}o����;�ľ�CJ��YY!��K�,>�&W�jժ�$K�2@�i�W�`榣�[?����I�S��`÷j��ù��­�D(B�W�p+�l8�z$-xཉ��c��}��/(�g����cl��'��r��d��ɡ	�1f�N�u;� ����y��o�*��aT��l���W�L�XΖ�Ӫ+�]_�ފDj���2�cs-Jq����=T�]m�̓&KN���1��������Jr�3�azQ}���PD����Տj�@#�j�}Q�C�p9-��QQ7�rQ����Xr�߅d����N�(����m(u�[�Ax|c��	kt�F 7�MҰ�i�9�0�{��aJ�Gm~��-��4t�Z�"���`;� �m�ؿ���͵ƒm�(�a���p"p�	�d�_�;iل'Y�:�ǟmα�G*�\ ��HE���pu�]u�s:h�����tl���Cm2!e�Ä�n$gnj��ts�J^�������p������D.�ٞ�^Q>
�\R�M(.߾��a��Q�c'�R�'�����+RO�f1+Ht�*����
"�E��Z�
P
E��|n�$�5����qH���t\���(�����A��RK9=+ ��{�=�����/��w�a�}C��N�bfSr�&g#�̬������i�7l���mN~u-;�;*�p�-�_�	�v���?�BS���y�hϴ�YV1��ͯ:�y���	��f���-�;d�H���P,J�B}�U-)Cm�LG�{q_�V-��V���	I�F�Y�q6����2��o�D۹W�D���z���'�6Y;�Z
!YjkY#!qq�0"�J��Ƚ���9��R])%�N�p��_�ԉY9�Ϗ���[;<#tS�=�4SW��-�2yT#W�=�"%����6Eh0l(R�U����a����<�8�����nN\g#���d1A��&:�3YG�����J�X(���BE�ޒ�$�$����F@h�^̈LA�K�@ʒf١��T��)���W/��,7a�.��z�y��^�*7��ݹ��͙���� `��wLZ���h