XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����E��4pC�rުN]��S�xyư�o)�WH��]���C��#�Q���/�%V��W���,?��qڽ��ǀM|��w��I��'P4�6� �_儸�,�;ɨ�|X��
�S�8��L���WsG�/~��2r��&s/q��@��lD�����'�X�	g��~��5�x�e�3����8��y]M{k��H�?� txn�E�}�s���b���"gҰ ��I�H������SO�Lh&���B���q��wg<}Q�!�7�e�㬿�i�\��K#N���������2<u��a�M��\��V�\:��V���É�l#x5�tNތp�aT�-���ԑ�N?bh��@-�W�*b�3a�	�!�䏄��,�]a�c�IV�b=�����sf;�����t�)���Fc ���!Us��al��^:(���V�[����$Y�0rh�4?yݙ��>��YLPǧO��`�����"n{�A�z��|A�-�$��s�}��|T�˼kSa��&��g�h�(ؽB:Bˈ�2�E�>�WG��v����X�`�}��Ů�#��KG��_*N$0��:}��uf�14��G�,�����.z8�+�>��`��Oe��v�3��f�;����0�@K4/Y�`��$��M`{���H �)4��������h�l32�:������������8�.�{�@�����N6	��(ڽ��'$�3}׮�V�OSK�91�L��)��C��:�z�.�3>�M�]��XlxVHYEB    28ae     b60����5���s(�$c^��+HL�YyY���d�u��BW^&�,�B0G�<�︘��h7� �\ �J{����ϲ�>,�#$8x�9!�*���P�`Bt쎽�DO���b�m44E�>f�Ÿ�X����b�Ga��<G��E噖�"�\���}�s��໋�X���"v��s�C"AJi�U7"�[d2���x��@��R��K#X0(
�t�;Q����4·���#Y95|��	�&�S��ϞO�ꂂ��T��4N�juZ��*����Qβ�-�i	w�
\~�C�k�zK��K��D���',�D��	�@Dq���$ؔk7S�������ͮ@$�W��\rw�?�Q��%3�"���I$�:k��pu�z-�sVS6R��}�N��� Hi⊺��;FW:T��v.؆9d�������� �0B���
t�SD�8My����R�h�V���J2�x{�"d�v�Ǉ��Y�t(B��	��k���iX��|<3*�L[��q|�7�/ʧH��Lb�5�mAkHK��1nq��Pn���+C�k����w�����S���E�qHxUAc$N�[*�����]{����o��6q��`2��(�1�meH/3'_c-v�(Ӊc<򗧑LNd�/������f��uIB�����8>���ԙg��P���{hw�0�Rs8��'��tdI����{����&��r��|3������$�6b�k�WRso��Zj�␀�ф
��.ӧ9��Ĥ�1�v����^|Ӵ�:>E:����T�b�j��*�@QP�{�zr0<�N���mm Y�d�}��Q��&�u��M�/P��`�uEGO��՜�Ӱ�dn�ύK)���8>3��QA	��T�%�D��� ��J4�}Q�C�Fg{ ��w���~}lQ҂�~�������#.};��x<�Ýn`����i�W?5t��c4��j�o��t�P�ދ����2�e�X8xs�̛�������X;$����s�:�o�`�Gsş)������nYT�2�zs��m�g�$BaI�X��k˻�O(�/n�r�W�3�8��#>*��W.y��_3�DN$����	\�p3��W�z�$��p��<Z*!�'[�7�]�J����+�<�y�WT|Dӌ�!@־
�βءҍ6� 脬=�<�M�ɇk^ʌW��� m�|���*��ߚڂ���v�FeA>�:�+&N�i���A`���9��#�.��/�ȩ����yU��fPJ��@Z~�A�:O���y�l
�AFq��	��n�Z6M��}&b,��!�
�W%l��Y
��5%�~-tN�o�u�_�#�OF��q�ԉ�^h(����0�Wf7�}���CϖW���۟��E����n�FRʶ���{	�GX}|̽`4,W۪/k�}��
tg�k�Q���F0�:�biuf@`�?9r���X�g��r�����K�]��O[;ø����q��VNӮ���x(5�)���RR��i�C���hp%aඏ/�z�612��-�K�?,�n�kG�V���#<p}����G�"A-]�y��Ք���E_�=�N7g��}B����&�؋�Q5����'�0(�o�*���7�-Ϟ"��Z�+��:� W��Q��h �,Pgȇ�AP���y[m�b����9Ǥ��W���jG@��׎�,�����ʪ;3{���k2,-��/��<�7Z_<��c�1��Ƴ������p�i�Wfj@�N����Q���zP�S6�Y�K/g���w�"W�T��!�N�'Xu��E���C���O+l�HmX����A}�E�����o��лμ}xc��@)�Ѧ<YD�'�-�����`��
َB���-w �*,&���
�L�sS�6�����<0�$���ʐ�d!i���8,�(�����׏^�7ڴAK/f�ҝ�����ج�7�8���1v�r@�!�E��*.b��W�'௉%H;��?���~���k��DUp��Ǔ�U�_�-�(��W������eYeA1��o�) WG��ڴt@ 5�sw5�Y����&��텹�M����u][�C��V�h�!0�wr��ƪiaD�+�#�2W���������X���ֵ���w#~��VIAү2��T�p	j��a0V괏>�1S�N��\���g��d!����R	�Ii�=��7.���B(�3`���=���s�rhl!F`E'G��J���Q�m��D��PB#t��I���Eu)��[�:� �|m��P�pN�-��K]��)!���fp1e���@Գ�Tf5��]mL/���Z!�Sr�@x���DK���g��#�׀�i]�ΉU�_W�TPY6 �0�aq�l�P"�Cʻ/C��)U-1QQ1V6ԝbqs�Ԣޅo�`EQ���e��M�:<��Y�|�ؘ�5��wt+���]�"��,u�O<��gޭ	��M�0��r�X{`��>\��Pl�??�6IƎ=�2l֟���4)�c�3�"��05�ރ����f�,�F�(6�O��Y<�N}J���p=�zK�wI�όLu�%����Cc�#�ʏS��<IZ����%�S���,|0}#m��]N��`��E^�"8�[�l��Yj�a��R���{ce��W�7�4
�0(�ؼu��Dú���^���Y����%����L�9���Z~���a���[���F�"i��*�3z'�e�D2�ͱ>��BX>N����e�}O������%�h~�`��"(�������g�A��Z֑Go������B+(T�x4H4������k0�Cɉ���0�����}j?�D������ ��Rп��췭z.H��xc$�^4Ԯ��!d�AL��