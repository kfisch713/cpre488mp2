XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����M����gȏ2��mu[�*���p<!2������x\*�̝���&��>�]/!��K��^hwO�L�dL��e�w�ض�p��@l�#�R�(RLi���r�/������8A�fw�Y��7ӎ�8ՙ��~#zĶd��,=�OQ�ש-\�5+�Ldow����ϢڮK�ՙW={M��	A��QG9}po1	����R(��������Co�>N	t}t�ιe��Z[���<�䜊ӵ\��Ið�)�(D|&+q�����s�¥����㳈Z�r��v鹁kABB�XB����9��Y�V�6#�a@_�K,�E'I���.�|�|�j�薀O��ԏ�����9�Ǽt!`�ι��3i�����4<��:lF|�:ѕ�~F}�o:�i�����\�)����bS,|�I_�=� NVT�(x6>0���y��z��Gs$u]���qՕZ�P�j:HC_����1�R{����;��*T�+|�о��o�~pQr	b����5�LB�l,s�� �����W�|GtF�VÌ'uDbk�i9n>��⒠Z.X�R�ʚx�l99�����[䠄q�f!'��r*Iu���M`�F�o�v�L�G7丱'k
��p*�h�����/��ҵ'��6�`>�~��ɉ|��A��G����nгBTs�%�̠_�:9�����=P� K�����w�>�D�HɪB�S�^u�+m}KRm��c���!�\q�60�,|�߲t`h�-��XlxVHYEB    39de    1170��yl��˾<9���R�ݭ�\�lBس�2_%U�bZ�9���k�rޟ�)�5Tfd{e�j��o��ZK��H���d=��iCq��m,��鋠ڐ���OE(��	��{k�C��e�?�K���b)������(���J��.!Pi)k���� �6Xm�������GMp�%�i;MF[a�m# �(�pnO�Z$�C%?��`1H?�y��¥�Eυ����s,?�>��$��w�4*��2>���-B݋	��R	��#>������p�kj&��R�3>>��&=��=qH���^x(t��"[���_��O^EMI�(�B*����Fд�����b�GX�6 3��2(��e�=�i1�I&A_|�@/��c���[���d`3�X����Ij����Y~&�B?B������֭��	��tu��5\���5
����"K?;�8?!���E�Ԭ���/����>J*�\a�vҝ�ӧp���n�#h�}�Gǯ)���C�Q�*������b�-�ll���p�%v������SSɦ*ަ��:�wݳk�Oo�o��`���'�&��v�[�g��u�x���U)�&NP5U���q�,��߂t�����u��O^M)q�4��#�H��>w�����~R`��&{��X��l�@u������7>��i��Q9��8��F���>���!��)�ݸ������ً�����b�}�Gݽ`�� ̫f	�(�
��e�����CTC���{��e��$nI.� �qv��ۉ%b粆�*�{A���gx;��@���r&���B�����0)���c�Iއ�y���1�hʅ���z<$N�g��s��Δ*Y�"9ªE���~%�5,�w��.���zQ��<o�`H��9��HMJ�I�"���ɔ`��糤��4����ͭ#�=+��]]Z��G։3�I����?!���;�u�l��&����h[yn�Ma��`����%��ۓ���NlÞ��#8����(Z<��>�2��� 2�hZ))gၙL	@�m�Yn��zq�k����w׎��٢_�U,�&4R�����Y������u�w�ES�H�${�I��0`.�r�(����mV��N+�ԙ)y(�u	P�J�#��� �	"� �:'�K=�u"�򴧲ߚ�>�/�ʲ���n������a�P[OH8K������l�P��5Z�<ȑ��}z��0z�V���[Y�M�/��f��t;8�0k�Z��Z[�=Кy%0�>
�T+c}��E.h�nsC�Y/�Ml�B�0�IT�ؗZ��^k�
<]���:�|̦�T#i�V��?S���	B��u���u@+�ڼ�XĚ��sӦ�ăn��(�Ww۔�-��\v_�SWw��OD��v��	��?���kt��7W\	i�`9�D���j��I>Dň��a�`e�"�����=-@�O��v�jn ��W72�S���� r+s�F� �KտB��� BB����prY%y�G�[z x������qŪ=����ĸ��j���|�Y�wMzbȇ��en4BK�x s����mE�6����]�t;�`2zԜ���+�.+�2g�$� |W1��o7��#����W�^^�S�5>O�t>���^����4������U{).WE����^��{�?�nO�ʰX���`=y�#>!FW`?�T�f��������f�j�Y/�Ygq���c��>����~����Ï) >����f��˫�1O8'O��)���g�w�����/VH�'#�Vcړsx��! �f�w���"����;�X��.'c#P�s.hh
�ϯ�'��C�YLҍ����)JIH���6~P���:�9�1����׳�a�����j%:N�#��}������2m����B�D8p��Y�wN�#�!U�dG��F=fV�P%1Z�.ٻ�sϾ� '��ޥ�F��Ѐh���K'"7�0 ��h�i��%�O�k#�5����>��Bjyo
a1;���M�'3�l�n����	 V�d��U��#�I��NS��Tǀ$�n0���SO:S�#����eY(iN�����C���a=�7B^J�V�K�ClwI2����%u=Y�jbJ�r�1ܶ,{nŽ�ɜk�����ą�:����x�)�(�0�7�y������7��m㋯���k�q��ِJBB֕���Y;���F��JC�B��\1mV��,ViM�6I��\j��&�s�c����_&NuC��1��,#�͐/�y�I&N_�Dq��㽣I�U��}r9@�f�z���	ɘw��H�*|����)��W|V��O !��O���PTE� �������a�̔�>=��s�A����7��I�� ��?�5���mr�5��s�XD�:o���z�̊l��O�ԓ�#��(x)v���x%��\fA6�ӂBq���;F�d��-�
���9�B�(9N��S�
�_��ת��L�JPK�#M�;Wu2�㟀lvu�4�V�W!5�C�#�P����$�]�����������,�(��HŐ
c���d��;��<��z¶L���]>��yM�����mIbMH[G�*y��Ϛ2����=���Ĳ��-㰮#�����v;���]]�PdOB��ᰏÇ�V��RZz�,F�KY�P^Y��펛���S�W�Z�﯐I8�lNa,BH�䟬9._B!{_���a�H�m)�ӑ`�(ߥ�w"��ٕ��D>��H��j���ASr��8�O&c�mt��O� ��?�t����6�rK�Jj!�0"v���G~�i/��F;@^B6�G�"�R�v�ZwYy!R ����9U�s���@�Z�)�Ћ�U/Q��/�C�Ć����k%x����.Rʻ��R��Oj�ˇc���Vxu�Z�2-6��P�a���t��C�1i�w���'AP�ty�Yj��W>�}� z�)���n��Nߘ���m�8.K�=T|p���UQ4o�A;�fҬ�q�Ly��:�����&T;��Z���;gU]���Q7�ݽ������!3���R�ˉpei,�g�����L�U��ڕ�BS��b��ך�1�K��ҁrF����f<�g��(�������'��{+U��.�߱a�
�:��:�ǀە��`랠:�o���d�ɀG�#�ͫڐ�E���������W��s��u�20I��&�Co��.Y�"h{�5E���觑#r��ž������^[r�Q��A�?��n�bζ'����Ep�,=J� l��6�*H�$5$��p����𧨔�3e�������w茗���%�����μ\ �hU� ���ڡ�΂f�ʼ�=�$�LAAJeuj����������3��`��p�n�
�)�<��^ف��J�w�r�;��ޛ!7l��ݓ޾�q��wH�F�-����T�a�"�9č��
 F�>03j
J:���`�~<�="kJ@�@F�B��;�&�IP�T���5��$c��3�,s����E���v��u���t��� )��ij�1���[����y{��0Zt�U����rQR��Md�c��
2u��x����DoO��Z��.�=���FM���h2n0q�gſ۳�Ҧ�h(�/�'�M�ਥ�D���s�,#g��і��I'/x;t��<f��������,&�nk\$WL��̼��m����D-��a�PC�v�l�bM!�8�0��͠�hV�C\��>Wq�`n�>�0�"D���A� ��h�C����\��U�G�~���Wm�ŧS0Vɪ�'�nҼ�E��v�@�`v�d��="��4`���"Z:��� !i��\|Y$SɝY7��M����~׳�ы��Gf]�̡(���ص�n;A��5�R�K�&	*j��������������|L�%�������"��f֣ ��[�1mu������y��ՙ���~$�����	Ӛ	�c���YT׼ypb��l�"~���Ȟ����qn��W���/P[M��F�Gq��A֏Е[r���j9���h��(�����9�yC�4�^�VO*Pt����hi��P���Mvri6�E�b����,�i�h�.�T^�a��E����;%c ����d�7"o\[wm�1ݢ��N���_�G��[��c���^�˰�0S
�)֤�x��r��;���i���jx�2S���r���Ǎ:�n���Yw���b��>�F��x:��~���9-���=XcY\��,d%�f�6@9�C������|���D��S-��T��^ɗ)�<�Lw��22�7Ǻ��U$�Y�.�S�PD\c�"�Ok�y�x��w(�� p�x2��k��!㧒ь��a<� ��r�K�/�/��:Yj��