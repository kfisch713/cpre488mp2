XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~t�[^��x�!5��0d ��,s�<��1P��s葡 M�_�u��������0}�//쳤^� �L�A2mP�1��W82{0W�e�YTX]AJm�ZS,X��3)�􁿇 C5yQ}W�jn�pGt�=6�ǡř23e<dW���L�꩓���ܪ�z�����QN��i�CXѼ��*(+ ��
�m�X��l��r#��jLǤOd�Ց��a�NO�JAl|ϨC�����9�.o�N�1.����@$>s[{rS�a�?��b���H�i����4�ѭ^���R�KB��i��dz�	]��%d�����
^$-�]A0{D�W��|��6��=����B��3���~��Ud�,��֞$��W�:�g���!��Tu�bu<є]0����+�W�?O� ���R�*��Q������ցR&Ri֨���=��D��Nmb�7~ЅK:��;2=�қ��sg����=�� �}��}�y��2�/ڵ)�oֱ�_���ӭ����N�앆���s\~�S�ټS,�d_YĴ���,J:�[��W=��7��v��N�"Ǯ��r�yoo�8�B4��P��k|�	�U�Hhh���P5�}ҌL�����1H}O�Y`o�P���8r`L7Z�M�'��c���į���i):m�Ғ=��T���# �@
D7UW9�;'>�ʰ �hO��WN�o_vg�}�� C���6�g�5�,���l^IX��dX݃k`mK�O��1��X�.[}�vCNW��&j��GL�M��XlxVHYEB    1448     800Wڌ��pz{*K�Y�����i���Åy�&j���Q+�ݪڊ6s�g=z���c�<��P�W��Ntq��d�����^f�&ȼ����ID��P��5䁜�=M�{�]]�0�DY(��}���T�A5���*`5K>���cq9����y�+R��n�1�g��ѿ�g��St�2�?V��m)�歺�� jӳ1��p�SڐlG������L[:|y@<��R�Êm��Ϛ+̠1}��vf��j�zpk$���|O)a$��@�����-�/�c~�윪#���*c3)}�B�2�U���⮏�f��@,�0��?�f�q]�"RU CY ���.R:�xQi��#vu}^r��%�9ܘ9�w�&�% ������Ya�\���F�D>���jR.3�t�chP��ѻ��{wi^��b��ߖ�d��������?�"���8�����a��WtG%Q:�b! 6/NQ�qQ��-*sGb���8Ʉ�n�U���ɝH��I���b�sn��&p^�&7���d��Qk�D�Q�S��_̼��ҫ�r�bH%��x��j�Ϸڱc��ω!�U�ݨ�7��(����·Z./񂯜�\բ�[�q	u�J���v�\�&Ȝ�@ʂ}�T��t�tC����~vv�2�r��	~@�	?68o������A��8x���=�Z�QK��F�+�M�����`�@-�=Ե�zh̴����.�V	�'��ӽ ��-���k�L%U�Xtk���v �~�BRz�p�R;&l]���էd �9�$��>7��R�L-_):8�MНm)��yb;7�_���Z��7Ն���X�Y,-�/���)~Uk�**�E�U�pE�Bc}?xAմ��� fG�1��a2�>�.����A���/g�}%��Xԓl^�^ �A��D��pe�$J`t-ns1) ��O����.B���ƥ�mC��b� \����U;��F�r{���Leusќ"�	 �DRr�O��ҷ(���']2͟H`➋6��	���R@���I�k�{W)'�%��z{K�=��V��p��yV-���GlT��%'i��>L_���A-TmM5h�'�f�n����R-�ء��)=���ηB�g��=dZl��|3�f
� ����%��S�G�v�ِAZ��Q�q��g��CQ�l'�	���.����~X
@P�	�e�q�|c��df�(����^������QI'�Ș {�n��hd����|�\5z�w��q#��#�-�:�IW����+�|Vg`���J��~�d���T=Q���Ar6��c�jqԠ���`�΁�*4��ǺTK0\jRD����{-��2YE𣛞��N�V!t�ݎ�!f�E�� b��r�O��ڔ>�iqf�	Qa���c�~��w�x�B��cP����Evg8�,�7���=��]^Q��O6i�L��<��4fkV����f	GXw�S���e6�T�}4�6Q��B9`�@��t)v��n�74����9�mX]�ԏsI�k�*w7Q��$��1���̪�{����uX�� :Wm���}L�5���b�{��[�� '����Ξ��������I▲ٟ8�7���#�j^�����V�^>��
�*�����pȞy�p�x���8�pߏ=�c���`l}�W�H�q�$vR�@53�Z9�� ��U3%�әC�5�'f�i�J�:�Skн��k�?��n�C�.���@
I8��p�=�f:+�آ(�����PAϩ쯍Ī���i��`.�*�?�xwĥs�y례=ݴ�B�y!�x��Ǝ8i1�����m5� xr���^�or���eu@Ղ������'���j�B꒷]$'�%`�i�G�;r�=���4�4{p��<�J)�س�zs�\��{�1�4jol{z��*���A�핳
'��>	�wW���.�ǔ�]x�oߐ�8,��O7���U�V���MW$�<<e/�9�J�E��f%.���ᙏ�¿�g