XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(+��d_h�J3`������n�'D��#u�H��}�6������u"�b���x i-?ao)D����6�U!�{�YH60C���sD?�����0#���s�����s�3����tg������Į-M��E�|;��L� ��%P9�!�����`�;�_�����A�M��r�W�V.���*I��g'��\�f@�Ir�
i.��LSb@��<߻'0Q�[�Y�bi��^���z��X�S��:��HjE��b��q�gj)D	s���|RlK^H��v�h:+?�3a%ڴ)��ײ�>�Bh�z�":�H��F+�B/��|j�L���{��'��{�*Q� fХ3K�1J�@QT��aꁎf96�S��WT���c�w�P�`K��k$��Zmޑ����*}dRᓷ�p�v���}���EYR�r@��L:VN�]�'��/�!����?����v���Ǘ-�Z+�Sξ�r�����(nsA`ޓ��B���'�G~L��RxS.<c���t��Q�T��x*;�ߌMˏ��rr#�g� ��T��/ϝ�9�L�M`fړj?<.�.Za�r�Y����x��f��%瘟#2�6��P��Y�'�_1L+" ^�k�fh���GjdRMYM���D".Y}��y���s�ƭ?���Y�e8O.T'��"�$�a
���!� ���0L�r�jo����a����v��M�(3m$�{���
k��t�`�u��|^vw��:�9 ��@�-�%�NS\�����טh�S��AXlxVHYEB    1ea4     920Т%�}�n:_��
����s\U(�����������x�g��x��w:c���h	̔���{TQ�����t@g{���7c�P��������~��Ł�gw}oɈz���)%EEl�P������'�[�3�d{�b����8z�ջP6_siY�5�"���c�Vtn�W��Ȍ���z�ku��7T�|��4��[@-��]�K�����1l���ξ�$�p�Y�Y�:w�ib�CC	�뷛E9'~[�.\�S�u�@&�:C�=>~kw)>VPh�#��Iz�Nm�W������N3KJOr#���?>F3@��w�p�6?��^w��Щ�	�6No�M]�t|��8���ޜ،��h���iZ)�=��Z���񫾪��Ck�E�Jhƫ�u�f{S4n�)�3nC��]��'�	ۂ��l��7��"=�	`)�37J�x6��^����
�����0�&�QC̪���\a'�֤ ��f���ϫ�	0p��������J�I�Z�a�Q5U�v3�y�փ�aW�N�ƾ��;#r��P<T�-͒Yf�s�Q꥙L��@K��T�V�CU-���.d�b'Z��l��,b��%_�����X?y��*=���e`��VF&� �H>�*a�h|�s}��--S2��޸me�4y�p�O7�Ol�N�}�-N����!-})�w��m�������o���Fև��z��>\�꠰mә/ù�|�d'���h)r���:9���2!�t
Oy���}䢛�b��A��<lXZ��^���"q�ңV��)���T7`��[�y�-�����K	�s]�<i�6r�ش���$ɞ��^��A�Rފ�1�n���v����7�l/m�T_��^�]�Aj���}�V�L��-��A'�J��ba���D��V�U�j.�aʋ~��ޢ����l�@�-�+���Dƞn�x��.��� �9x],Kh�c`]K$Z(NWv|+ܣ@�G���dg'ܿ#"���q�H�����rT��6g֧M�������&w``�+����ښ�W�����q`+6,w��@sM���3����^"�O�bcm?T{~][8Ws�n�0�6"��Ə1)V��}��������!�('�ץ�{P��qH9Ǟ8��~LG�f������95EcӔ���\�(Zh6���I�7G�4�/J�A���Ḑ5�M���٭a3BT���9��k��Ŧ�j�����<8���6=�Kt.��c7�t$��M��00x�΃K���	ݹ\�[f����>ͫN�Ө���N���ve�W�Θ�Gs�E1,Q9(��#���y:,�|�;G���7����zMq���=��h� ��&�kG�q`HW9s�r��sF��(�D�����"�M��(R�*Y�/�@F=�E_��ix-L�~5�������Ea=���|�0���٧#rୀ�
9����@m�ɍ�SPB=6Վ��Kꃧ��^����ѡ��-=K��K`Gk2�e�f���.�����vnf���ٹ3O���9N̒�Mb�t�ߧ]o�����8�]"�E{k����Q�y�yG`g�Ը&D_�d�H$K�I����)�����j+������
�l��=�@�S67�0�a���m�o�2Zs�������+�{	���#-���m�kaW�m���l�@��D�5������~r�!o�Vү���@ݼA��{J���� 8I5��$�� �>(�I$��Ju���^��o�����FnD��8�%W2�	�ߡ�.x(��ȝ9�JAߎ4c$a����1�n|����l��V·A��칉��6M5��an��U���ݳ(�� И$��ݣ��̥�\ș'�[w�h���*0U*�5y��HPK@���BXlz�	/wb�'���!h?��D�\���5�O �	�\u�%��3
=�XF^�J���2-Fo��&^:t��
dJ�9���1b�U����4��Z�~��	g5�cF�}��fWq���+�AQ�4%<��h�x,��.ԧ�o)�n��X����������M�w�87R�Y4�CԢ��k�h�l��Hx��F0�D1: T�k�����5_���<?x�i�m��^u�4x�%�}�>bor� 3��Z��5�NU���L웻�15�C���W�s|HG���/���}��7I5�@j"
� ��	u�m�:�X3��f�Wr��g�9�lE���IH2���1��Q>��N/������il`K�@�т��ۼ��X�������y�����GȔe!���Z���~hRi�����rf�t�n��o%��ܴD�