XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w�#�i�4�.S���\=X���� ��ZTآٞ�n��`lL�nM��~]f4q�,6Ďl�s�ó@����lVTߋ~����)���>��ȩ�2�E�0s�h���TaѠ�6ƔPa��/�F��qH�n���i��giʚbBF�����}CJ�밾W>�����֗LI�VFgY�Ι?��P}�~���BMx�3TՏ�G88.�<��K�MGtA(]�����˧N��8���&T��-��Sj~�����o:����sDb7���e�r��B��l������
;�� �Υ�	J-�CZ<S�qg�(��}��QB`��qgFX=F+dJ4�!�)˘�]T��B��Ξ�`(�#�p/�f���'/)/
1��Ȱ�5�h*'5�O�yWz>���
�z�k7�Tdl�u���9��	�Pj��M������T�3����z��w�����i�!�4��xu/�]͚QlܮR^��?��F��d8��ULQ�����Q��aR~h�(�o.�1��.����uf1��~��_�������� O���>��|nS��n�w���-� �յ!��T5ԁ��!t��'��0K��q�#�P+H[��`Ca��8��F��'�H$
��0:��~v��>���T��捴p
��i[��[}:ө�.<�d��(�~Dh�/�B�ƺ��FWS�n9A���7ˡ)�u�Lxpo�\K��I���Ω��f�0�%��O'���ɓ$]4�d�XlxVHYEB    95d3    18d0ei+����Г\��� _B�@��wu�;F��P�WG�YB�h[�'.y�d�����~	������:��7}@]S���,�M����N��ܷkqC�T��^�����B�h�:6!�K"������܅y�դ�W�q&��8"�Et?j������7x��s�x@@Vk�Q`�A�n���;����!Df��(�5�U��T�7�vT���%�@�ƾ�<��;�%��g�l5Hԃ���k��¢�1�����EI*��q�ҭE��}N"���#�f���	`� ��xK(6dh�2��O(i��vN�;+��cR�#��e��*3�6��4�r��(:�3c�n��q��o:����K�Z�.��%_�O�7@���1{�xh\F:� � nebq��Y+�������5��6rF����.`\�S!�����&�*$���h����l�=>���BU�Nm���ܺ�t��(�}�0.v�֒�&\Fө,���{�Mdt9ڶ�3��c�;��?L�C��+�C�j�w�E�H+*���p�ߪ��OP.n��h�(;f�% �pvH;�]	!��mݣo���xr`� �;@�V�ܧ��ԋ��ɇ/����X��V)���g;��jc���T����X�[Y��{�+c�*���ft�a�ƪ�a�����_��<(��3�G�da$/�_#]�d���iۿZ{YMF�E��S�p��MRӲ�v�3�K2����,�vq� �1Sm�SV=�S��f9�F���~���+yix��Z��t���Rߊ!I��Av�Wí��<�Ai�z���	��T�[i�I�f�	4�u��P��WJ�k���c�/�>2ی��=��\�y�R��]-d�e��e���>���E���d�}?��*u���IgYeuH	<�}ɥ������	�v�=�镨A��w�����1�&6ܚ��𰘗��S��,��H��U��G���v5��Ȳ��9�w�M�����G������d���7P�詻Ӛg���Ė��qo�ck�7�j/v�{K�v�uKn���x6M������!��@�������p�"/EÒ~�:(����`TZ�CJsTzs?kYę��=�CsW���qf'sa5��8�y<j*v(�s)T�= ��<�K�%����M��uA��2,� ��56hџ�-�.^k���o 7ɣ'-E[M�1��Uo��`�J��a��Xcݍ=�T����M��d��w+�=
΢Z\-��'̙�~V#&�@��pfk�i*Ǚr�f�x_N;���Ck+\f�M��]!20� ~z�J.��@c�[�[��US�@$���0����厤�䉐���#E�sϋz�v�ϙ����+Yp׆���]ez���9gi4v�}��F����ӷkY�D_]2�~6�'��:#��M��ңm���M�������g�c�r������"!H~��|�*���q������������/�Nsɟ {$ ���1,�Zb<�8_��Y<���wIC�m��"�/�`�"/�,���3ǵ��G�GA֚x8�z�Z�)��xAf�ϑ���xp&^�<������S�T��৷gD���̩�Y�]M�
Aw&� (���Wa�o���u��D�G�EH�S6���s��w1�Ll����0ġ]��yjM�ț�L:�#vz�E�g�ú㍻��i9W��w"^�&��%�^ b�ۭCK��aB��<��C2��*�]%��V��xC�j��˳}�L3�R��O������W��	���}��s{p���FC�mЯ�k��ϝ�����x��s�x��_�o+j��h�iV*}�_q9OO
l�9�� o7�i���)`{�JL�wA��d3��T�"�����1&J3(ۥ�ZU�O���F��,(�����:/�	�� �����9��,��cz��ε@�\7y��@�$��,�]?����k�V�K��;w��F�v�."{np���z�1(,��׮����]-�pF�:�*ߝV孅�nM�n5Jo�J��m�t]r�B%��'�
�u��MQ���LQT5�x	�����KmY�t��:�g�p��;��:���C�`.�8�l�:�lA�3�$ք�C!?m�w�yo��t��xy�<�3�q���ؒ�Ű��ەX�JZ[�H�F{3ܶtrO�����]�4(DT��C�)T�G�~M�F������j�/�~���5Pu��vMF]k�'WLZ�mf	�%M7~�F�ߐ�Y�3Ս�����Qzx�j m���<XU���$Q������V.<)�w�ܺ_yR&ڽ�J੔�H��~�&�� k߆�{I�1QQ�1*�U�w_�צH<V�>]���s���j��E�X�I���4%I����$���!��37y{�-C&�7A���BG�XZ��
uD���I�a�B�j�U�|�2��Wŷ����K֐k.�{�j�'��U����XL��
�{�fקE�(����r�'��W*��$#q[�J�B��Y8rB���x�<�~�x���ޅf*��^^��@O���"hIg��.K��:�
Z��R���膱��`S���g5ש3]:�� �_�����#�} ��5�2"/?���q5����u��h%|X�L�ܴn�n]ݶ���`�d��m�[���V�_�ľKa� $����eR�L��_Z���kk��H��Գqwz�?d��b����r��)��s�5Jkh�[@����7o5FdnHhq$3yÃ��xD�*��N�+�����Y��-*j��S�n�=���-[�e����R�������iC�Մ����DF�
y^�b�\PW�S~���DQ�wd�|�.#nh�lj���8��Z�����.�.n���W�6�d�{/��[;gu{"��޹Ql9_:
�����]4��;��8���Ri!$ Z�2����x9d�"~b���?�?�]��R��6nk���6e&� �A����z��>�Dmo��>f�:��.* o�Hz�$���n���������c�ߪp�����ܓ�I
T��߅F����2�a_k'-��}��">�Փ�$�G����k����IqW2��$��T�G@^rjY��Y���6TQP�? ��R���h ��3R5�HU��D�=��f�	A�ZA# �����H�V�|�{k%� ��G֔z��Ǿ��,�2�S�pp�K�)���UU���׫��"gP-U��������,��#e&�X�Y�?@�TV�T۠�^��v¶�
ah���,1��0pS��arTpu+FqY����D��jg�?�q;:��^0K�uT�{�k3[�|�*�>ʶ��R!��t�bo��${�-i�� oz�R.����VS^�T
���W���$�)�����ƒ'$Rl��!|Zn�8]8�i��-�H�2 ��ʇZ.7V�h�d�y���t��b�da'������0�����0�"v��L���ۀM�,�d䁕~,M��}�<v�p���\E�A��+ ��⢲�[*(ғE.��ᨩ�f�+�ӝ@��zHl�(��#&�h#�dOAO��DZK��۝B�F�7"{�B�B��R����˲��3? �rÈ���硬�7%�$l/�0�o
G9�y~/�w�P�ѫX�c5��o<�����s�ؖs9E|�zn�=��`�Y�VK�&rL4ps{����9���_/������`I�[5��6��4�c�8Ľբ�I�o�&�0�z��'���O�W�;�f?<Ex� øB��,��>G�5��ѻ�1>�������tOo�8_�[�I2�(���p�9����H��*�V�gW}R���(���K,�ĜLt��߷Ū�}cvY� I:vt�<WF4�Α;��\m�4g_��H�r�@���}OI��:�0�Ql�����R!�#�D�4q��F]NIP]H.�\�ɜ�l���',�|�mX���p2��,�¯���i�,k�@r�b��\��0W/�"G�H����'����w�BV���>>���׭8��8������t�	l)=T5�5����iG_ss�3G�=� f��7���>�+��s����H?EH�����ڳˍ����Xe�-[� OtnM�Oh�g��rd0~pҹ3�UC� ayͅ���W����	�XS�V��8���0���z��*��2�.�J�4�v\�!��Ql҆E�w�7ȕpq_��Ur�����i�	kY3�F��LP�����4[(�r1�#�$�������� �aƜQ7���
��T2�vF���<	_�ۑ3�a��#|f��_���ĻBBbm���w}O��i��	�$@#t=#����s�6�W�\��VL�;i�ɉ��Z	��Bη�$��>|���Y������ ;�^ɢ���1i?�ԗ�z\e��RT��#��S'+�XڳY�Vu�1?�g��G��V�x��O�%� �T+C�]	V߳���ʒ�����x:����3;Jw���'ݯ������ׂ��N��ɯ�I��G�&<���������M���O�[���8�X��5�Hv��öŗ�a����,���&��=��s��M�c3�k��G�M��i |�q%Q����(���!���M�u��W�oq��#�
���0dY+�6vI�	�ܔ�'�	�B��?�%���TBfZ7��X܉}�z��]���K�|'��Q_�5�Lb�_,r�D���m�d��e�Q`R���u$�w`�n�tmri�8��i�pM>o�2�rM�3tO�և��bg�O�1׹'�!��g�:�{qP ��J�mZ��j�L�7�Ŷ��Eݙq�K�zGV��u=?:[�`?p:���i�k�z�̢d� �|40��aK2��N"�o���R���S0��j�䜊MG����Aٌ8���V���~r��V �w)O)�˽K��6Cu�Y���Mo�|�wB�@����3|*�HS��{��k� 
�d&τ��w]���N����딨�&ͬj.�+O�g���H��"R.7��{��Ų�
=	�OɟBq�NF{�!4���XٰO6�*���!�jJ�׮JT��d˴���<�ҴyJ��M7����V�;#5/£�y4������J ����� �SE>�<s�Z�.�K�`��(�0�Q�'Ig���$�j(�������H�꩛����(����R��C��"�Eu�a}v��6�X�=��!���NP����a��X�ΠR�:[��NI�b��8dXe\��#��P�\1���b, "�!U�W[I���~���,,~����#`��uʹI���܏!�쏡	��Q�L�Ae�ؗ1�7�A�s'���VJ�e��ߩ��f�#��2�����S;0]�����!t�Q��[�z7]�5�'�FQ����>�H�Eן�oկ����YU���T<'v��cBT�Y�{'?���V��Uv�Sj`�f��H� ��j^Jræ���~eq8߉2�������d\-~��1����\�v�kT���EJbK$/v�*��+ejoɟ�+侊�v���^�0�$��A%RL�`.�X�2�rE��Α�l��1�fC3阃��{��"G���Ϸ�v�D� �r��������B�r:���rwL�!��,ϼ4������Ѭ�>/�GZ�#=DH/6���E+�{K��}�xN1fa�:��b"c^:đ��R^�#7�,�mhk�m�d�m��s�C�I}v����4���ڈ�����3�8&�40�D�h�6���Q����%�b}�Ҕ��Go-�px��4e��/pQŦٲ~/j�o������/��������vE7�=D��V���:�I�`��d���������@�[���@c�{?k�t����w!�����Z�#`)}n��'�Ʌ|e��q=�Ƕ��?+Lno4���� |��v�2����_w�*��	{K�d��\n�nS�//�3.&�pG���[�#��1^��>��<��J��?��i��!���K�a�;�u�eT�e*�ܖ!}S����eyu�o ���Q�6�J&�޼����,��^x(�eQ��g�G��a}ܛ��C�(�Ċ�Q<�V�%m���I�Ͻ8��(՟�m�^1�af����� 1,� Ƹ����v�2B\^j�5�� 1[�6����#[��񾮠�ݐ�I�?��g���h�2���ءr��}���ex����9������&)�����r���<�?*�^��o	dc<�^��螇�n)�KO��m꒭��m���a�m(��hbvE�M�=�Y���Ki�D�B�d
�	�