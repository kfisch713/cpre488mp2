XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e���"�bދ�Z�y$N�2lp������8I�Ӹ�M`�d�[c��PSS-6�sX|'�b �{@���ϦVv��|��S�ǐ �Y�����Y���/�}����N����ueV_�������z��MP���Gt��2PI��P[�yb�P�P���j�X��8c��{{��A٘����2�k�4B'��ա|v���q/C��C�\;�CpQD�[�# ��}���U� �84M��K��p
M���s[�fv�Y-��ƈ3 ��]�yl)�Nk1�������2H�0���R^î#��Y'�2��_�`˃�����o�V�8P�O�c���?�N�UB�!2�� j�����Kcg��<�W�s�6����:��V$�a�S��i��k0L@��ǌ��7�bm�g�נO�۲�=��N�V� ,�B����u/#9�{ |pN�'4��/k!�+�o�|����"��>��(���K2�Vo�������L!�Ji��������eݪA��7�ԃ���ջ/�g�5�z��PP��h�BĨz��NA�1��(�X�4��D����3�Y�'�������T�y��b�!H�f�ԣ��z� *G�,�d�	���Ơ�T�o��&"}a_#J�yټ�p)J^bE=N�&�����)It�qb(Ϊaۊ�"R���oҹ��n� "Jo)��=�2/����������"�k,"�R�*��/I
H�����Ӆ���BD��Ѥ�1x���0XlxVHYEB    2b75     cd0��6�i����Ǽh���r%������;�ѕ���9��~T��T�e �5�Rl9 �.U�m�"�WQe�Ғ%�d��Z�+H��6D����B�,Ot���q�~����7E����.ׂ�H<�M�^V�9����q�'��
Dc��i�q�d�Cƪ*�@�GE�:TI�$~�zbIU����_s�/K�I��t�b��:=Hh��-�W�,�	jW�� �p�	j(p�1f'�U��K9�E2���`����K"�(�ߒK"���{{�h=�������.�7}��i+��f��_E)��l@,�����s#�UD*��ۆ�>�U�?t.kr12���1�Xa�h����]87q�:$x�Ƈ�5���<�ĕi,���*�Fi,��6Bg�6�*�$�{���J�*`�6��=B�VO��`N��jT k��n�s�1E\�aRU_e�
���p2�@���s�D>Ɯ��\0�m�O��&��٧a���se"�>|�T}�s8��y�W]7���&���V<Vd5���IE?�F�0�$ܨ��E� �I�ձ'V�5k���sE��5:�����IK�r��L��%���U�K�6A�����C܉f��{_p�ͤ�q�nd2�v�-��>Nu�T�{q��)�e��"%�_~ȊdOP��$��^��*|Fsr�����w�'��Wb��_]̱�Y,%�
�MBk߁�!?�b>�Ž4I���F_r�S�V�%�^�2(�̦�w��Wf�u�='s*�{�~�j�u� �S��Wl�E�ƺ�rV]���XS�&h���c��d���XY����n����s\j�9^u� Z�� ��Z^׺O`�\,�4�_���7�/�K�(�Z�|�8�i�&����)v���7��g#��1\=�)�Z��j���2�I�]U����y��&G��`ń7��JS�~�B���&��l5?�$���:��:�݀{2��-
a�#	W�S��գ	��a���Ne�xH��E����h��07�^p��,�����-�_���@�����䆡\���V��D��K}�2i�J�/Zk�6�A���l�gʁ������vn�&�TDZ�\��$�)5 � �/���M^ ����,ik$ �����z%
r���e�������+��$�
鐓ļ;>��)YGo2���O Am��x��Y=���S�=�ş`gg.�wï��ù C�E�u�b�/�'���<OLG�^=Ͼ+�l��9)���;�U�m$:dR+�)�i����$��0�U�ۘ@�	�w6љ�Y�,:<�y��G>����m�����믴�P*�`�`.[[ *�c�ô�y3"o=`3���%���4�������P�ik���2(9�:�4�MO��l=��{ڠ����*�[�f��H������؃a���3~1?�ee�&�l[K�]<���d��zs�zp|	_���5q�{ۡ]���$���������`M�F�����c=����G;G��=����f�蔭]L����U���gR��C���:8���ˠ����i�$S���J9"�T��r=oAhz�}�9�m��\X�ёD���u����Tf��-U�5����4�0�5u/�!c[C�C�sH;��g����$~F�,ds��$�s�	�m�qzI��u��88l{1�UdB��Cm��
sŁ��a#�o�!w�2d����rR���82G��z���Z젮Z���.�3lLd��0����'�Ń��;X�������;�	<I\2TwjG1�+�چD��O��mJ�a�y"C�AEޔ��}hc~��Q�W��>~ž�0�X�^�v������Fn�M������L����㓹&��xz�� ��,��[�����,G�&@�My���O��E�V���+��p`���I�lJ�"��B�f�E�1�����QHv+�v�<?kkkO� ?0��)d��zFr���>��)�Hc��O�0�l���A��R&,<�G���ྉ���wl�y�"Ač�2U*��|:*��Ԡ͓�Lu��/շ���K��4-�A݊"��Ť��n\9�c�	1��e����ANp�ME��Ű�!_Y�D�g�sJ���
IG��b����bU`���Y��fb�o��K�(X8;��K�Ro���"da�Bs����D��~�!�2a�IW������E�g��95�ȁ�\��>���y#� #oh��L��e�įа� �U�!4\˲�Y3�|k7�H4��c�Іb$�Z�1@Kt��LEe�!�/U����SO���{�H�/��S�2�2BlZsj������n��S���9���̷����M0,a�.Al2"����*S2�U˖"I)i����KU|>_�'�@_��ן�a��	rR�\�ƾCbV�	���RƔ���X"�)c���?�FM�N��F^g|t!~��mSA�s.���l-S"�C��.6����)S&q�������F�%S:��JWw�:��?�IN�
M�r|�=���:�Z5J�\WB8�f�q����SՅo��k_`�}|��J
����ʇ�j�;8�:r��p�}�&Ur�����vή���*�����@Y�yU�N���9<=�FE��[,c�_Xr�N��Ş��.�0���ݲ�n�鹵��q)]��:�B� F�,�e�g���� �7iW���FW˼7��V��;���9~LXk� �-�,�n�47����5U4v�<��,� ��"��M+v���QV�ؚ���iE���'�m|(����� 9:�Fޖ/f�ѕ�ޟ5"v�׫H������Qr1\��d�ՅSIo���h�ݲƑ���DD�RH�U�ͼގǜ�!�m��� ezф?�?YJ0���U������LT����w^���0в?���%�R�}��wܮ~�9����|Wr���S�¿��%ɦ�S�L���p�}��3=h:ͷ���;4A؛�x��%< �P�a���%#�55m�ژ�MO$mh�Ml�OE ��h��('��μs7�faQX���x졳��۪��,�s�,�.{:���a���پ��<� �����|�6�Gn���+o�J�E���O�BE,�k{¢` FI�'_g*#�[�Tڦu�XPy�qDGA���4n�����V����bo�V�4l�e?1V�_�[�S3&G�R��J��7e�)<C����,
lXCČ��VZ��m��P�Q�7y�^�;_����\[�َ�\9�6