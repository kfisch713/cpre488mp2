XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b�T������Pa�Ft��uȟ�N��يlxJ2Ж���E�?�y/�]V��R���.x��@2d�=���|�8�� ����(쐬-�|yշhv�0�N�X�W�Aq�fU��\L�U����mw.�\��Np���a<�+	4���yD��C]}~���j��{
�Z|":̾�Mt���BG��66Wܨz $$[z��w�0S���VN�U�q{h��x�/�(%�<����-Tۊ��&{?�"�]
��C�W���.%P���vHW�Hi��4�	iq���t�0V�SցJ�Ho�l�(��	�s�2�;��ԇ����,������7�^��C�?�yJ��� A;�io��k0
ᶾ���(̿XX|!�L�E�5�fe&�-,e$,�f�4�'3����+
����}%n�[�_j!O����X	I�/iS)M@h����t�!=�
�Z<���{�+_�t���wu]�6����f6�څ�dX'/,`�@�DGʶ��ї�^��
z�ic]a#���И��4Z��h��6�}�vd��|6bB�Zp����I~��f#�{��s�g��gf��g�h�S%D�:��1����n��{ƀױFl�k���m�֐Sٶ5t}C�Ό7��[P��|�N%E��0���M8Z��r���L�qa���'��o�gjC ����j �����>�5���)V���Ӫ+̄�f���	Q�D�5�,6c>�g������&H�}}+�e�Iip-#(��XQ��x1(�e
	�-8�,eU�>�XlxVHYEB     f9d     6c0ͩ�g�uPx)����=�͙2+7��Q&p����V�kSǟ�ֽ����e �����=�ӊs8�˻�lh�0.`��*���WiF!��8��qF[����n�0��<��< �����M[���2Δ�m
Bd�� ;#��H�s�Ξ�`>6�l�C-<�s@�р"qpl��K�:�,�O���&GJ�M	U�+�A�"�
���Ɉ6���91+~'§|�R�V�f�4qv5^g�,uV��˞z󣅭��f^gs/SM�m"9�Btퟆr��b�w�4�)�������+2uv e+���\x>Gĳ�WѫA�y7�+���Y�������r6������p n�?�}��@�i®I�}wNx����]F$��C��� �3^���iϦh�,e^f�T2\T�d��'��hH�tu�"�AM�g��℘������C��g��8ɐMO��V+��l܃� >��Ի)�C;y5��v��/��I;�"�	i
2^��t��2�'�#6��� �3PmP�7�,��#\��8�o/]�/ ���7���;�>G���8����j��D4(A�69���1�-hlmEM�������({��u��s_�I1�@���MCEa��ǡI;�^�T��_ZC�Z����W�=�'ث�F��d�9Sb��)M�ĉRL,���.۵�}�8�ߡR�$��\�T�����y��/j;�|� ۳|�?�����!�*b<�Fgq�4�@Dhv�JC�����q��Q�pͭ/�k���#����¨�}S{8�[]�A'�eK��;��8�B�n��Y������cz�'~2��������D��wg��p�}�֞���g�a#;����#�dߖ�G�e�OK�;6�M#E��tL��+#ԘC��(%c�<��ay�,��2����T'��K��W�T��Z>�.�@|���vި �&2��:ϻʧhŽ�^�����/y��0�o���<64�޷�P_��0x=���FpC��|�Q�I�<���΂	�
/�{���%Rs��ׄ�\�x��@I��Ñ+�Es�'���5h''0�2�����y���z?%�^)n�9����ܰIc)���5��%Smi�`B:���1'���좻ތ
?�wd"j���-�A�W<c�L,K�����Ӵ�|���]��YԦ�������-��,jM2Qƞ����������F]l{u�1���{7[Ϣ���B���^ۗ�O
�|،�
�}G5���&�㢣F�9H|Q)�4-���ĺ��\�26��c��S�2���z}� *).w�5$�[��	�� 8��L��"uM:�[ja:�����<�ϗr�n#XqfѾ_�N�J�b')l��6'6MV�JFd�G$�t]�����J�5�:��wB����F��>�����M�P�qէ3Q
|ѕ��S�?���|}�����y�7�gS�F{��6�5��B�U��ɟ��9R�6�\j�~ɒ�����X��(,:I��@��b�ؒ�H��Sw�c�9��oHNA����/MO� 3��\�a����&�(j�B�f�����i�1�?���BHTʿ)����.ր�vxT�}��s��^|�ظ�8�D�Dg~����t� y�i�s�l�F�0���@�y���jDĳ��ް�#x�#@R`�}(�T�,˓TF���m�4.��BPa���