XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/z�۸7)�*F8J��b#!%`�A��5�lUܠǋ�Ұ�֑����`�f�劢�P�����L�ȫ� (���F9�N���jc�%/���� <����д o�ԎyC4����\�S]���x��h�U�6]��P�bƛ��tI[���h�(��d5��}�0�=���/�����o�IV=?� ���ENi�߂�d-����D�=��:[����v���%f�������A��iU�9� �d�."���"&B�k���z&(&�η��IU�G�G1A��p.xj��V?��ǧ�)�i�2jʝee8��;�`�_��{?��� ���T�^J=���K�
J9�<`f DW��ޖ�+�:��uW�}���4[���JS���MV�c���aD�b%z���{�:hE��o����c�;M
I����^��B��]s��XX��p</������g�k���>$ذ'\Ie�<L��^J2�1��4��W�;l96��X�Zs�<z��6��a�i�keY��MTObE)�a�w�a?�'b�ෝ�l��95%�׮߉w�1k��%�?���oq�źk�dg��1�C��m����>{7,�G6:ph�t��{.�a�G�J�)�u$n3T��`"���Ky��]�Q��"�jݓ�0��24�tvdӞ�2�ݢ���C)�_IE����p���lWU��S���<ޑ�����;`���<PiGb�:�|�r;�Դ#���!t�S)�}��;���XlxVHYEB    9fc7    1fd0�5��Ӿ����ǋ�}��㏿{~̓>�F9SC/�lf����E;qx�>i�*��^�Ӑәc��? ��'��`c���F�aD�
�3ҭ��H�[h7�@��瘈f�<��E��U����e�H�Ԟl� Tp��8�q�C�r����ۅA�j��Qܪ�����N#�/k��֔u��p�v�~��^�ֶ����O�k�D����Ϳ
����O�gH�@� .��s?"�8c�(u'Ԡ4� ���r�Y~�j0�>f��1�fE��,���ο�4L�����a��pX� ��L�݈�e	��۲�D3b�,�;X%�6^XҢ�*n�ZR��=b�-�!����u7\=0�I����-��w�ԹA��ى��hX��X2��-�'!���2z�����˘Y
��ܽ"�AI�¡;����a�����tRW�ˆ����,	��P>�x�n�<P	ʁ2�����i+ea0��m#2_1������|�r��D�֋��LBf����W������I[�VY����8?M�g���9V"���X�*���/,�8KU>#��t�;��\L��3 ���d�)2'������8�AnTƠ�@;3	�T+U�	)�~����7р�]�,�-+�f)�*!Vy�bF���T�%D��Øn��3�	�r�����>��p9a�
�MTcu@!�X|k�{��\tB�#�v�>,ZX�%��c���&�ks�3�6�؋df��E[��4�MKf+��8�?�*2����%�&�I���}L�r�,��� Z���Yl�${�X��1��dBk�/)R�@�L��8�v�����N�֬�eBލ��yXV*g�e���nP�T@�'�}�ю�J��A7��+"�՛u���G����&��y�1��ベ��s����-�)�d�z쮂����=I�\p��:%���ow��&�� PD�g0z� �����eT��o���3H�f�a}TW�Z���'̫��PNs�����-"�"����!�B0ɢ��'��W�q4�Mp�镤��ʟ	l���{�R��/��.7�^�K�d�ꀬ��TXZ��;��]�\�Y4����y����}%Zo����x!�|����9�|5H%R��ƽ�y::y5�Y�Y�L�-��� �H��49����ʏ[��
QN��reU�ۥ�^8�x��� �v:����%��A���`�/{,�!`Q��E�W�+����T7Է�����ᛲ+�����,\%B̭?��<7�G���t8p�Na���]�g9j;3l	�Q������S��>]�|ڞ��/�F�4u[�����_+�%�CQ1M�a�_�StjJi���˾m�f�m�=
_v�J.����M��WD뀰��=�x.\��Ƞ�`����OI~O�P#�s�d�!d��^����c[N�vB�W�k�n�>Ҡ�D\�L$����*r���hGgֆDDo�J`U��u���3��6���nL`n�� ���/��$C'��b6�O9絠X�����O(��(9Y{攀����Έ;�t0�(r�Jj�1���dJz7S��T+ƽ��Ey�wYv���A�3�s)������lM�H�%S�T��cqKf�P��[��S�A�#�y�D�Ok&"����a�	�k7Ç��9��P�`?�R�=Km Cq8J8��;J�6���a�־LHD2'�f�=}qg������0�D�6\�: %?Ԅ����QXj}��qz|�u�`^�-QAXf��{p6��Ӫ�:�
\G��t�[9+�w�����LO��L�V'�[�ƮN��,OuKVF�6�L��,=��7m���)m�Տρ�p"��Ei��ాS>`���x�ͽ+����ǒ/P��UǨ��xrG����� �[-!��x��lBФ�O�� ���������&�����&�yc��nr)K��	�ǜ%�ڪ.���>�f������F՚�`��YU�/��jb�߂ў|�o���6�'p�S ��s]�����Z�����15̖�7�7����lX�[;V�q��g}��D���$O����p#���g�'\�5QY���/n�_�3y�޴<"Xۈ����g�hS�[�6����U�G��_������G���
%S+J��S0�iroa.�v	@:�c��0B��T{�`u��re��^$�-k�̀ݡ�(+R���ו{��x�I��1��ό�5_�^,m��=��8.a�v��+���L#�jHÜJ�H9�Aȫ$g�YѨ�#*�T�SE�UPuĺ���*�0��S@\U[��0�ٱ.h5͈I�9H�t��H,T���t(�/<�(�,ZOU��^�m�]���X�� N�'hDI'ʯ���C�>P	_��n��o'���ɉ�)|���%��a���?��'BX���a#��x�%�v�/��("6�\�.��[ƛ�{��;r��ֲ/3�����>k�0k�����h|>!���}<�8#1i�p���=���5e�*ܒq�|"i��LB���%4��02p��N�GB�a�GĄM�ߛ���J��x���m�>ݝ\g���@���h�y�����W�W/f>�������1��Ғ|:�$�U�Ure� 0�ъ�_�2�*X�$�,e�8΢��=U�x���ۼ~F��m�#d���y�[��alo�-.�Y���Q�3�s�-�!���k�5Ay=ƸMZc���l����ĉоΗN����K��80��pg�#�:5��/@��7��\�7_=Y�	x�
αP<��dNؖ�2�V��d����/� �k�S��U�̥�7���\@&�Ѥ ���$��͹<m��w��ߨ��?�Ԯ�/�Sf��� Q����[7���_�O��#i�8#4Iq3��Y�e�)̍q9�=���'� 
��f�V�B�X�7:����?�̜A�s,r�
w�0$$��A�; mU�F�q1gNY��/�+�#Q�B��D��f��D���^����U
���/#�g�9�Z["��H�PA�V0�}�.A;>�BJw�o�8�(�s	���}���U�cۅ��$P��zͧו�����a��k-���
U$�}�l(�K&��h� ��Ҵ�)ϯ���#��~S��C���dB�Tg�օ���z��ǔ7��Z�-/�����	�㬱�>�|�=��۱��p#]�1Y����l���%��⃇=��Γ ˝���q����ф�����6X@Z���i vE��Z�r~�C�yV��q���,����7]�%l�l�୙�>�W\0L����I��6e��f�#�§]�G@�p!��pu��?»���d�3e� ,�Kf��K�W�)��x6��i:~�K��nr}�en59���}ވ"�2��~7��=wn�hǑ
��gd�$�],�B��j>Y��\��8ʜ���� g����q���Xy�;<[�k8�A-���h����M��d�8h	Z#�ߘ��׺����k;�>��o)Kߦ��f��)���j���l�s�|2��n`y�6����S�ZyO�)�ͯ
����m�e\'BU+Ec��#��P���U*��1]���
Q�L(��G��Y�8b��G@�Q�u�6§��2R�?�x��A���\\6?M��9�>�~|h�{3J��)�l3ʔ�puG���P)��:Ck��9X��o�I��AhQ��R>����rI�b�;/	%#5?�}=��:El���ΞEȯ��G�s�T���9Mc��܀������D�>��;}�jZ+�S�O�×fYs��)2G�lR���=�G@+��?'����냚�x�2���8�>�g�B�ɫNj�י�_ɟ�=�I�u�D^�Z����h����T�:�w@,p�&��-;��t�J�s�|���y%l�'�.x?8ۢ����n'����q�,h�^��L �����{���d� �튢:�
/SA��Z��;H� �a������["�;����TNa�&���_�*�s�l%��ʺP�h���2:���V6G��bꆶ�i@�	��4��	����k���U��ݛ]�h��k(%��7����Ά��M��n#��1-���`� $�_�s�����Y>C��ֹ�JX?�`����c2��w���@K����V%q-ï�O����_˛��|;� �	�{��]��?���}q��N��nz��L��xţ��ٯ�S�W,��c��۹h��}V��<��>8��xl�+~e2}E�^�2��P)E��[�z���m;J�9Ruݥ�/�+ee.�jba�HD�q²�U���L���[���sLG��l��ja���R�������ww,�ň��U4M�DwC��4��� W�y�EEx�tTynqP��ln��A����~��
�-��U���u�ԇ�jRT@s�������\����~Y�ߟ���Bd�pomRA�;�,��K���mty&�%����oS_�m.�zSv��l�}+����Eד���6��V�]���i�/��lB�BiM���3����U��׸�β7���v�?�-x������ԇ1^�]�qȜuF�)�Cr� �P��kg/9lN�������O�ɌcYUA�FM�=�w{c���zO��2�a���J�Yn�{�Bκ��B��&�}_� o� 'L��M7\�u��f�V5�QZ<���Ů�acjP�G^ʍȔ�Wgm+��ki�zoq������^�!5�[��m��7�|V�T��Ene(^%p}�s�^�;O�m��QB6Q�Դa`�/��t���x�f*��U+Yf�ڴ�y�� ���,C�� cx�V�)�hH��G1�l`ye��r�Y`#��(:��%�H)�dF����Q,�*�)��W���͈�mO�ᐺg�^̃G�D�|iɚL��GY�m��:pY=M預�
�-��xǁ?�1u����T&P�8a��>��1_}��}_B�� <=�N����
N����(��}���(�I�)5�p��5�皯t��*�L_��)�줈yJ�h���K#�v��������LHx?���Y\��j~��v��b����C�|лW]'���/��<o����5X撓������]8
m@u�.��Ğ�Ѩ����eŎ�ˣ�f��:g�ml��E�@�l�,x����k�6�����D(�,�8�|��L��Q�Z���@bΒdT�!��v ���;��Nh$���]AK�>C? ����FQ���xq���A�H�ww��C�H��)�#B�X��APw����`@��E8��<�-i5����
(�{��kW���#
�Km�w��K�^�]���]�Ұ3
����+�������)��:C�4�ូ��Qk_�l8�P�nT�2�"<TfJ<�K�Z���������0�<�/�s�s�n��n��?k{��k���A �Ec���~��Yb�2wKx6O,�@Њr�_X�J�x�o��οmd�__C1�u�7�#ň�Y����l<����E�V"���C{b���C��t���O^�4����_،�T�^YB�)	�H��b�]c�e��q�K��	@[�x�a�vOc�=ә�|>�N�e=�� �B.�`3��x@<�S���[t�qc��"���fc��cl |���ܔ�4__]'xD�ߢ��djаm��Ėw_0$�Ð��G�"%}-�#�C\�fӿ�p�[���?_6���Qvz�+h����?iY�.,b
8�q�&(ֈ�p�:�d$IQ��
~�Q�3��zcP��R`)��Y�н�36�`���Yk2]�^&|�,�|�_5gT��l��q���B���)p�As+��X�2���(�Ӷ�*gU����ϛ�Ǫ*��h�~��N��	3�Ch���0:ɯѧM��D=�`�~9��$x b�^P�M|ZМ"�Cp�A�Mņ�����(V��nX���Y���6Ƹ����.J� o>%Aq��f5f��Mb�<�*��\j�aъ+����3����P�^Ͳ	���{0�[��:��+x���q)�7�3R���@"/'���zv��2�l�y2��M��O�G�� BX��������*�:?N��]��vq��1��/H}!�ى���~`���w%��yD�:��^��"<���9*�{�svě�5�r�y�g��ک#Xz���Kԟ��4����N�\�4)�d
y��Xj�8��\"�	�`���Ʊ�G�j�!K��J5�`_0��n�}8����>��Źޚ�{ZO��:�"tw�yT�R�#�Y�J'��ŵ+�D�^���_��5�>�^+(�
���|�<
V��;��1>7WH��'8��ҸE���"�yn��N���yJT�Ag�'��qZ��I��}���iP�W��h�CZ�+���ҙp�x�]ja_�����<B����>x�^|���˱����R/��`�K���Ԕ�Ly3%e�MٶE�jɤ�B�D\�����`�.��8����@�C��U�K@,�o��b��}7x��d����������x�P��т�⪻�$�f�Z������Y�����Pehi{;5oYs��ږW�F����<<�K-��D���4�vF�vxiW� ���E�hoJ�:��k���(x��c�Y��w'�B,�Q�PX�,��r� �K2�#���F^�M?h��LOu6�HibD��T��ȹ3 Dc�f�n���һ5���(Đ#n�b�	�Nӳd�n �KI6oU8
�z-,(��zOc����ZZD�+\�O�9��'�"��jb�
������3iU���<��NEy�+�{w� �䔮FO�bZ-Ā���" �5	�쯽��:IK���+�1">x."��!��F�}�m�N����ϴ�̿	���'d�	�|��c�8��_׸�cW�-�K%JY�Mg�9.�'V+�l�v��1v�'$���EkʕEX.��u���:#Q���A�P�9ػ���,@�����g�d���'g͢8E��*JJ�������,�Sl{{�p(~�I�.	��P*��!���[ڱ�RL��EK��Z���8��qѭt��`,��@G���AL�5�X��=��7E#�If󮗿k-ޚN��Ň��yiҲ���wΤ?�@���Rs��+��s�V��1��8���B���~�Z���-��\be���%����2�{������}ɲ�:������?��9���Qrv���?Ӫ@M�@��gi̜��c��Ҿ �F�h�X��k����#�mn�u�>?ȷ��l`��G��$�G�KIq��2Un�9N�:'c�qZVr���x�Y1x���G�����tY�-3�o��]0x�&�:']4�d���V`�f�ݗ~aW[�E�^hX}�۷�|�0��ի@As*pI�tPg��.~�O�W�Y�#G�1w ��^�h�p9�>�}�P�X�=��^TޢK�����:N��>��M!��`�3��~�:ԔB��e��bBG.��H>ڗ7%̥�=H{ƃc"���5����^=���/	i�4�T���F˻I�+^C��ig���y��<��ڐ2Q�[X-��	������^gsO�Mk�iev�߻M�B�Ԓ���ƀ6��F����_�ז_�Z���#h�^G	<��V(����$���b1�S=�U��_�Z����"R�����H��gnF��X�p6�۷5n����2+bJtQ�X���l�_Tt����i��|O5N��� seA3���Z8)r
��^!5������3&h� ���y��b[��ڤ����l��������'u��t�Z�,Ӥ�P���Xї�d{&�~ ����,��]�.����Q_n�&y��Zu��p���m	���QG�]X&.���l����`�ie@m�rl" ��;����۽K��\��Z> Sσ��z=j��b��̞Qؽ �X��nJg�]E�!!'Q�G5?`���W!
��a���������+[���R�-��z\�o�7�´ڈ�@$»�'\"\�#Gנ9�ʚf�P����U(�΂�ð�n�S�K�XܽA&<��l]5;i��5^�\�"����JU�