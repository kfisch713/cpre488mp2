XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����R�h� NX� �uo���Uz�,�
DbܔD��o�|�"N/�#�ᮽ&�݄4��W�;#��������4[͈A�_��tu[��ub��P�n@*h�b����KmP�dCɾ���׫�vyI��W�S��D9��)3Q�5ݞ�'��D6�*.���l<��|rTjl�rt$
���SLC�tC�y=��En/���i+w��~pFB�>)A�=��
&2�?�4WZ	X�3���g"ˬ�j���I��W�P��`<�#cy��9�PY]�_��p���hѱmw�:a�J�,<�������F��t*}��ԉ�2�����w?�2���.��'���q�Ũ'cH��f �`Tcr�A�������k�1�$�9b��S�=��=캻*F��.�7�zɞ�����θ�M�D#�O'����]%cc�:?}bQS9��S[�mu�Z�;�w!�Ǖ.ߜ���6*hB�boD�-�`���%b#�&2�mQ�_�Ff�@g�ﳔ��vIQ���+�h�H9�ӳ��W��ظ�Y�u�cM"/��ϭ-4��c���q��v��9Jrg�H�9!2�+U���p��,�v�{b������2`Ty���1�	�0�:�Ys��*:*J��>}��8�dK�w�#�c�����X�"Im*,F\MN���+S��cpG�]��U=`���*�)t!����_vY���t�Z2����E�9����L�e���ʲ9+9�	��ƕ}�]k���~�=�"��XlxVHYEB    6315    1790L0�%l�5*��Za�68�#�}9�9g@��8P^'��b�v�����Y��2�pz�+�O]�oct?��L�ݷ$Xw0��@β� Oj����/*Ww�ΣZd*���Ll5�U��?�d�J�a�����C��g�i�iv��M��W5L�Q�쪬j�*a�<R[�?�DBB�E6�p�E�\Q�Td��sm�2E�g8� N���.�E�*[���Q��M�O����fO�1�Jg#w�T�?��ˈH����;���v��D��eN�d��!;�S��[7ޚM*j`�F$�QX'B�Ǹg������
���5�sl{� q����Q]i/����/3�G�=NU�xn��O�e�K��;8m�%D+5裄�����$a��6А�1�F������_��VCgF$o���L�n^N��N��"ӳ��eZ&h��0Ŷ}ڝ���my���f��H`��N�@�?��G��?�i��l�tW��iFt�R�1V|
ɱ����$�K�w5Cq�|)L�ǋ�W�������s=����7�c!S�s���YѾ*'WO�ܵ�`9{��6zL�h�I7�:�*{߻�b�*�s�P��߿�Aw.��Zk��	:jV̮~���b�ï}�`����ᗥ�jS{�*�(g# �a�Ӿe�<n��·T�Y6�C�\��~��w��t�[cu�(�u�=TctPҢE`����P��q�l�:!y�l��c۷�Z3鑐#���텿S��� C6@l�>8�>D���Ӄj�ʔvl�X�Qw�����|� b�>�zcTWA	B\��fXh��o�e�6�B߯��b��{��v6�N�T��Vܭ�M�����eyU�$1�������
���T��2���_뼹z]�r"��6�p��&'�D�h�{ĝ��g���KԤ��<$���8�ڳ�d�s����)�qӇ?�˾G���TJZ4B$e�ϳ2z�湈ߴC5��v�d!��,�eJJzT�s~!˧��Z2-GT�;j���t8M����ݾxS���OC���)˶OIvW�ukuۗ`B�����(z��|0�8<�(�ix�,�5ߖ��J٬?�
B�_alF��/T&����P�j�ǹYpx��XE�p�&��3��w�](�S^�Lrhg�\*�0��P�>$���!{cc��'��������uWQY?(Q�k�GO*!6C�3%;��+���a��\�}��5e�x�X��\X�+�,���"�����6q��~dw>R���-��;
?&��/2ד��;6�������'6��A<��z5���8S�N���g�fe�� (��<���y��
v�]�����[�:�Y^A�?	m&�����{[#��^�i�42�ȓ6�_���?���ֈ���.b�*��=��_w�q|��BY���"}Z�^��냘������e ��	���qJ.�~1�'�S�����#.�覶N�^�����0<�B�@�����k�&��1G�@!�Z�tд���kn��@����f==�2ͮ��sk_`�U�F��V�Mh7N4��a�W�ծrU�(��%�R��<�#Җ�[ X.���E#$��$s�Sw��Fe������'��*��;XA�L���yg�8�h��n�	]
J+h�泔�(�W�좻�Fҿ��z�
���J*��Nkwy&��^�]O���{��eB
�Ml^WpGI ��9���s�_?��g��}t�n�>��g�Kwzy���.���Wc���s�pi��h\��`���*��ͣd�����w��W�=)d[Ey���1��/ݢP��f��3�WC��=�Mh��*�捁�f^�h�TS����[wZA��nz�{E��v!>��2�̓CE�-��i�;�)��y��f���J�[��yK�m�ǺZö��Q��f�W
	���	��g!���������l-���U��ı��G-���lgS�Ҳ����}K�9C� �2�;�'TW�ճ��mA��n(��	
	��Չ9k�0��*4,ڸq�s�`�5Mɯ�=��� ��o`R���#R��3 �����~�U*
����V��(����w6�����-4��ӫ@ EB7PU]fØ5F*�:kq�\�V*b"��SV쬌���L�C�����O&�%S�uzge�3}�Ny�����ܺ(��M��	[��=����^[TI���hT+[=|oS�J�+Eff�� �ߢ�E���\w�a6�8�z���n�O�	���� �$t�cd��m��`[S�/��LxTj��,�j0�{V��x'G�@N�d��e��4Kf6h���I���n����E��mҁ��.��Ҝ���Y6�Y���MVxܴ \���t芗�dWx�@}�h��R&��K�	o���
àꖁ+�'�y��8W߼+�5��s"�6�Y��<���!�T��y��#&  c!�Oƿ�}o��=I�FD���&�k=.3#U�bs--�7˼j���M��Wl�������l���#��U~/�BѪ���g�L�u�����4����g)`�����ޡZ���g`<(Cj��	�E��bك�mIo�۲�?6�͟�TZp�_n�8��odG�z�kh����ލ��G���e��W�9�{�͎��S�\ˬp�Ěj[�5�Ȇ`^3؅O��p{�0l�kޯv�E ]�+��5p�CC���3I�01��j�W���#���`0�� ��ў��F��b���/ s ��S��U2�����+`0H\��ش���$wD��T�����fN��hcB�!� �Ɋ�f�I0R�8��Cn�W��En=�ԺM����JY����,˘9P����ڂ����H�_y�R���M	y�m��S!3�ƈ!�iDt=��E1/�b4�%�/��}���P�{C�9aEH�겎s��?vU,:�^.�%AL,K�xőd�;�G�@����0yC~�
L���*a�[o������3��WPR�<X��>YyL�r$�*RM2U�,��|y��d��ij��_1p>��t���{�aY�x�:�� ?F�;�9�$�,E�#Ӯ��T=��k��`�t�Dp�fE�{�@���ݒ�#d�e9W�I���������΂��	����5�b����e���nDxw^�x=���n�d�B�k���G2 Ź!��P��0����Nyɬ������;l�3q��Ķ0F6]צ-�0�����b��?��+�i�q67�HY�º ���k%#T]:�n'�H�����c�%���x&�P�3������;���s��( {;/wEZ�^�nc��g�^��+�#=�".�Ď`�Ll��K�f%�R����(������2��k��c��N-4J��p+���E��v��TuyS�,�]~� 2b�)ߚ7�T�^!���UI�V�'��j�Hj�>�?���=�*Cs�w�g:
Z�*)�*���I��B@R�Cl����j�Įg�ZY%�R;��-��+��+:,'T�Tp��r��Ic˖Lr�8��iq�$��7|;6`��gb�*�Mo4=x.�b��,<�"�x�^`A:��Ufmϑ��, R*�"���v��֓W~����y�)U��v�6�#t�؎���4�˲��u�z����Y�l�*1�}l��h=jV�J�S��N�Z������NT�F�g'���.ۍ�f��J�*����Zʜ}-��Me}GZ�3v�ǲA�ͮ�m���A�'�||ڄ�L��¯�i�Br�7�3�aU�h��G����
���W���x5�8R�S}�P��"�p��e�?����wPS$���_��ߥa��9Fz�
��#�Hsu�x�I���`O�=x����X1A�
�D�b�t��y�1�X�l�\dy;#�����0'�*[�."ٺ��zۆ�8��VMs��\ۓ`�4#|t��M)�0`rkU��Ҡ��7�a�뽘Ua�8v��X��e� ��g���-���Q�Vm�����HC����`=�=��n?R�N����mp���2��0,G��d�ȷ����_믋v�ܰ�)���!-�ҥ�&S�
P�n�&�M�VW�I������^��;8� >Ey�ݪ(��d�ʴ���~ɒ���ȳ���^�C�qL����ԭ%&Oqza����Lq�i�LS-<�zjU�L�d�O�r�D~��C��ƕ\ne�9&�R]�� Ff��������uu7�ANx��5�)	A������Lf�)+ ��#1I���%���?p8^�����Yy�ѹc.�_�.�54���F�0�ք6��C�a�<�0;��p�e��fX�X�̈́��l�U�kC��G���F�c* +.�&�Y�~�eV��d��J�[Z�a�;?� a[u�U�@ˡ(��rmU��L���	��*� s��N�S�Bz�&>�=<��� ��!���P����b�H�h���U�O���9�{��Y�n�֌nsw�ڨ��uN[U*�om����-ɓt�En!X'w�L�Wg2)�l�
 K��������E����
ִ�| ��3Dd���7.ʁ���J���.LpC�O���
���\����yּ���A�����{�S��_��`����V��*��<�ǧ�3� Ҭ?ƒ�OMo��E1س�X��4Y��j��fz���?+G��G��]Q�W�#8><�%)L-��z�*8�,s}�"��L�0��5��Ao��'|�6E+�w#n�^#LF�n]5��ALh��#�����)X��_L�Y5��ױp���t;H#ЎD��$��Vіk4��<�i[���T��:|@�@9��vAe�"�E~h� -��͆[���4\�V?���� ��$M��̹��G�ˑ ����x�r͍^O3ށ��	�~�,�����|w*3{F&�,��Ԭ
"�#Ґ��P��%�ԫ��|_rڋ�}�+n)w�}~��:�	;s@�B�_��|�8��ͳ�$�f{h�=\��"E
]�W�fb�h;d��W�;R�$�Ag岕7/T�mM�;2mK���ԯe5F�5�|�<)�(����PM��HC<�����s(.���0�A���YԖ� �y�O����*`�/-�?Gs��`�D߾�)~ſ@I�4y0���CV�uɫ|�8��:�v�f{��*�c�kS��L\�.���.�:�W�҈�\{��
�K�dO�j���f��s̏��"����PE��]O�+��W�(�.��\.]�H-���a&��Y܎<�/1��{^f�y4x���P�s�s%\h��:0+�l-�l���!/�,ݟ:3�s�"3�D�[ai��ze*j2�eL��BG�*6`��f���}��W�9�)�u��B�ƥF�Xv��V�O8�;�k�q����ed�����}�f1 �-4녞�`��I�C�O�/>�,=�� ���-�mO�. qx�~��z��«���I��b�l/S��[H,�x�4g9��b��o��gÉkcn�H�6.AHi�P�i�l����N`xs���w����b��sZJ֦�"��I���?������#�l�Fh�dt? Z��A�]��焑ilqBN��qD4����qH���c�2A�ъ��m�u�Q%I1� 6��9��or�b��'��B���ܨ*�xJ��i8��ƞ�|����[,s_;g�}������~J�]RDV�g�Q�����ZA�� Y��9q��,�f�b��c��6,�6"�n&z�WB�ӓ���|.3�|*���iG�Z��ԩpDR*O�p�
?1�AX�'��XGA�W�9��L8�5IrP��/���l� [wX� ͗�Y�|�ƹdJ�;��V��
��-�m�*y�<��!�^_����ف�y�_��y�1��Q�?���`���\�u'h]r���\�1;���e��!t4ɘ� ��l�̗��ѹ��}�1��E3}�
q��Y�HboK87� aҗdP����U�