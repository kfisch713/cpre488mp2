XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��urۼ"դ΃@NgU&��VQmCܹ�g�a���	�E�&ۤJb�?���a6Lo��T
s_*� >ΕHl=>�U��<�"�ĹZ����i���������WS�90���8(Ën��i�N�0j�(�B���8�����DK~��x���8������˵$WL<�=���"{��_R!��(a^���ɖ�ĉ��x�[����!���*
�f֡���H5%�Н�Rg�⒟ ��͍��S�ߩZ"~0�o���r!��"�hPY�am�~.;��f��'P���)�.ڣMJ�RY	��(��e��Y���<�F��_z�#<���NL���E5*w}+���:ͳ0�A�-���Q\,Mtܛn�F,~̢�w��9�Dv ⷅ����2����Ih��H��]UC��ȗk�w��#)m"��]��U�.�J^�a�������1S���� i�W��M#���I�z�Sĩ���QI?a���W���Fixõ~Wc�]-h��������y�p%7��?��b`�$p]ٺݤ�M%�~]qķ�{�A�CL!�o�p�k�KJ@��md�*M$�;}M*o��eBKY��4)�Tf<f_Ug���iݞDyL��qW-܍`����q�%�xm9M3n#9���i�k�{t����-��Q��r
��3��&��l����e�Nr�Q�c�./�+��K�C�U)�v����'�_�#���o���Иc-�i�|Ny4��|����۽(X_"��9"��P����N�XlxVHYEB    1853     8104^�4�Ku�y�|�Q��q�.r��n�%����{8��
�f!-�U�/��Q��KC�ʢ���es^�x�1�o�l���0x�Bq����׶蹆s�<^���QO�A��yy�7��4�L�'.5a��������%M��&;;�7��l�7d�ޓ� w&�$�,w��X��B5#�U��lȞ���je�?�� 7�t$}�<�'�v�T��V��иKe���өx!$���幍�����/�+�b���>�0�x��RS�>��ϟ���U��xМ������7���IU�a����4�\�_���kc���N�=���h��{4��t�s�f���!*e&Ͼe��� �d�E�A(]�pA�!G&���Ng�Gۣ}�zĲ�->�P����h7ZDğ�jR��>$U��Zy�i�"킷��NЮ�N��
��1�$�i�,Wm��!�|F�6��>WAc�&��o�5���Rn�;3mm��e�����<F��_�<��T����P8��E�j4��z�7cG�]NY�yLB�ֳ�+ķ��Ε֚2L D^4�׌�C�J�r�T��1E�2�ao�p�,�8����e�-�y��,|��I2���Ǵ'~�Y��W��w��1z^��8SܫѴA{�#M���Ԭ7(�b�Y��G����&��7�����}e�u�p��Cud0�����T�)���E'����{G�J����J>�*�̗A�8�XL�i���"L�f<�&S���xmo�ZwE�1�ؓ�k@��6���<�����#XvwIkGz�6�nl$��!��4�0<��9H�Q�OzvM҂�b4cN1�1b�����S���DԢGx��+��+9�7�����7)%M�a�]n�;�m�>���c���n��c8? /8۳����P�cҢ�}��;5�Bi	������Eb��&�v���UV�@�u��댴 �/a8�2I�qk�Y`i�r{6��"b����$��s(�C8Ԉ�Tl�1m���9�4�x��"O��|���F}�D
��Ś"�N�i\��ʺ��ȵ ���v,SL�7V�&޷Iz�PO�A�,�+���ꗐ����MZ/~�}����9UR mCeK��#X���=�Xq�����	��]�n"a��^��l�if�2�.�����	c�m�Uv�n�/��.C^���_����a�ȸbC��Q5�F�������H��3	�u n`JF����D"̔_j���,Y�)�:��1:�w��#C��Eq��.���n����GZ�e8����(�;��'|�Q9{��vב���Q.�F�`���ĳ=�UX�.�lAl�a� �~q��F:9�km[�i�18&�(�<�L�(<$�¡з��*NA�[ N�g���Uu~���Ti���qF��!�h'ƙ5�ig�'�l�<�8EgV	1�'�ȱ�豚��L�l����[
E-S�5ɩ�M� �U+�RE��Po����΍�0Bm���4T5(��׿R�4Ʀ�<T͔z<\�ȩ�A�R��z�AO},�Si$�}���O[�V{�Y���M�ވ�.�4<U��7J�rn�o��e�HWL6J�:�'�j@)`��#�3T]��)G�QL����U�he����A^�;���q&��l:��9�-fz$9� ����9pR4ro����C��)�bJ&�b��|$��t%�>��m�b���
�FV//HR|t�А��Y}�&t����O��4�p���y���4��A��V���8�Be� ����c�'�	jB���C&��/0�FR`'�S�|�W�S���~b�ųw:�[�O����q21yV���#(I᳋�X��g����wk$��#ŷ)Ԑ�(I��ɛ�O0�R�|Q�R�[������ƾ4��N/oL��t���дշ_������oyG�'�<�|	~��4��ӄ��e�Q>�DJl�z,Y���Tm�b=$uW�d����,����,�'�pK4�%~����	��?��Ĥ	���"���oc�)�