XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,�1)(�<P�zĮ۾W�.ш�\H~ٍƅyI����M�Z���k-��v靝��|栣)��]��� �hp���>���������Z�V��j��C��f?�hG���>�
l4��Z�4k�����R;�W�˔�ޢ��"W�c�y2i\�~m��3��V����C7�����=�i~�������Q��\"��Ie�#OHGA��h���ŀ%ٙ�����k-~���_�;�X2�UЋMko�s��t��b�A������5�1
0����k�@��>�g#K�@z\נ�#�⋠��}M��H������A-t][��}�D�l@R�w¤nÛ��Go�C��� j�y�x���Sv�x��g�������)&T9�R�g��ȥ,�{ϧG\�p�A{1���@�[�k��&2;mxym�_�6�cl�tBd�J]	��rH^r�a�m#W���0W������,D��HKWjf������k�*'���,�+�'�T�+o�y=�
c���l����7�P��S�:5�>��.l�uQ6 lio�,��dG��ښt�����v��؉fa��ќ�~=�-�B}��T�����0*�]�x�A/l�zQ�vn$��r�\i:���G9�Gp��L��;�_Ķ�OY�eD�ᡆ����5w�"���PM���]Oy��%�h=A�5[�t,�����Ko��/kGY�Ĳ��|��ɗ�	ILh9B�_�. u���0�	X.�� Ժ��H䕗��XlxVHYEB     e07     680�""/I�{TY���*�t��w��qh�k\���s[���+�#�84hU弜6�}��`��L�jLx� v
=�P-��^'mʿF2�\Mb�� ����cc�Iһ�0�Oʷe��@(�������F���Z˾�����������H)cz ZD��qIx��cx��w��N���kC�e�dȕ5�P$2�<"�8�]N+����i!��BW���F�aK���(>Թ���5:���FE�l�pA�[�Z�o�N���l���/�V�d��~8/8!����+՛~�v�J~&?�1����E�;���n 4�������eQ]����+�%$R�Yo�S�hԇE�&�s��8u��W��黑�.shm�-Kt��2�KN�b�[���N#�_��+];��ȣ�΃���HOM�����:^�zW��]d�A� 4���|$�]e�/,4^�u>_�������x{�E��a'�^��)<��;�{M3.�����;#��-�_�a'��������$$n���6Cwޤ'܀�x'?6"g�:�V?�����@��)����h�����:��C�ƥ�x��]�3�>�?#���Pw~쁘6 Ot��N[y���nc�Z�;�qy�`Ic�����K%z����*�:�	I�5)�ꇦZ�-p��A0i�i2P�����Z>���U,7c*'��L���t����+�� �m�� ����`�*��WZ�X�i���.��,w������#l!㎘��r�(E�Kr�ۯ��0d�B=k~�����(�w:���$�KTd�
��"���F?���~��\!��i�y�$z�4�5��|db�����iX�peT�����8q~�` �`4���.��)�!�n���b��s����k��v����(��.v!���>�Xa�e���3J�E��T�܏� M;n�Z*0��l����Y$]�1�]�>R��<?��؝d�w�]���Sj�j�v!2{�bO�du�ƽ��m��v�zat鲄��m��w�Mv��n"<K�d�&TE�;�AI�n���]2"����������,ޏ^2BP�h���Y`a?U�d��[�n�
����`J�@D0<e��h�<a�R�2�2����5T�iB�4�P����:E��#&wk���J���v����.C$V����#�L�@�
@��qj�f���~FSb�}=I�咫k�b
;)�߾�#�<	L3|��]C�-ݙ��A�z�d~��~���m��f/��'���_K6��L���������s"�8;��s�˗�	ͣ�9�����tM�(ୋ�/,������2 ���=P'ٳ>@���A�o�8b:65�1r�w�v�g����Z�Pќ�d�%����j�V�j>�p�j~���	�B��
0�����,��
�Ea�8u�iF〝W^F<z���j�k�TF%�\F&�-x8��<<�a�a�.)�}<�ɁZ��C�	�fu��p��� ,��	A,����k��i��>�F�g/j��+�8;j��\/o��B��~
�]l7�@������!X+�5l�-�w�Zl���.�j
e}(9��|�ɸM*D�u��i��}u	՞W(���5 �?N��f�Job�P!���v1����'8I�8�