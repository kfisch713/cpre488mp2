XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����}u�0x@���0T�a}\(6��b����=6�t�͂��5����w*0c���N(�g-8�J��:���r��~�T;��8��Y�������w#8��윽?����#! y�U�i����IE���+�	�03u�����P��u��]�[�	+'�$]|�H�lk��E~��Di��@%��Ձc�`��6٠x';�t����5�С����j�l�X�%�Qta��LIAR���?±L�'����v�!�6�K�A�<��Yj�7(���ɈN�^��Z(�U'�B�*e*&���y���7���x�8���5�=n�fVæ����ǀ��<�y�W�Q��8�4�*���ڴ����)����i��jV�h#0�J���=t/Ԗ��G�����x��m�k��?�ĿR$ r��Vn�F��}@�)%��yA�I�^����K�>7�y!��p�`�\�����4�5
��a�v�/�;Qׄ�2��z �P�<�eӘ��:bvmƴ5���1Y�9&�x t{��k����Mk3��1$�/��:
	!�0��N��!sx�%F�dp�7w}Ǳ �Zٝ�kr�-ySP��V�G.�\v��?�?�[g g�@d�W�|���^�X��n�(����2��4��I~�48{6�DrjV��J����Uo0��خ�
kQr�1�x&f���*	L��ҼE	�9����ȱ�#I��ë�)� c�/�do���2����&ޢ��ASM/A�ڊ$l *�4XlxVHYEB    7265    1660��u�+�P�k�V]K�B<�B�8��S��&�@b8�O;�8؂�N+.p����GL?�@1�|?/�;�B�>.G긗V1�����^��=���� ]��ў��o� �+�rv ���M�3og�d_��ӂ#�����w��nMU#jl�xI�,����3�\,�J;q^�mNJ	���!��y�ֻ����>�L�O����~��`n���XX�c���Y��k� �q��js�?���OKDN_��ܞ~yܠ��
UC����O:ef�H,�%�.WeԦ��61���+��#��Qc���0	sްw鰘z�-���4��{�C�%ݷHh�,<��yz�!�K�\�y��;{ل��q`s	V�����$Ëp�j���y�;{Io��w�n� �u�:�\FI�������5K'DP@��Y�� l\�!Ｔ���΀ȩ�$�G]e�^����>�Ц��+xֱ��~�c-�����M/�Ԯ
�-� �P@��<��)	!m�\|���4��2��O�����QT���1����Za���L4���_�5�	W�R�:s�JY�T�>f�?+
��̊d��,��u��&�.�qa���=k������A{�%yڙ��*�B���*\ ~KO֗�0���o� JS�]+b�p����8�3���r�n���?X�5qf������*�M��=�p��c��y���]�D�G;�+�E�z���"y�U��<�|�tV���!.���8ֆ5�ң%<��l��(C�V���Q��d�}0\�;E���<���m��-�#�E�{1"��g?�>|�t���c
"���?�py\x�p��G������L%��c�J]�N!� w���i�ݢ��2c��t!���
�=��S9cv�Zތ_��m���>D[ךʨ˳��Ø��Rl�����Ŷ}>�M�v�i��*�'8���Iר����M��<0����9�p��@Fi�Ȳ��;���Ei,�]����:��m j���vDA9��N�<�K��Ų�q{9����]x��%���N*�::��{�\P�+�X����ޠ�Ѽh;d!êkt���9��3��Nq���k� 2>։��/�2������7g�e�{���R���h���e����}^^ѭߑ`����d��Z��~��/�n[��O-��=�8�V#�;4�� �݋���Rǽ' +]���'g�hb��}���!�Ma��3R�ŉ���\���w���6<�D��	�3�>�x�.�QOn�+�!�h����9��,��}�z&"R<���}�]ߘH�**�ǉ��8�9!(e��r �0 �Ѩ.��.����[HA��C�$&�S��o#���J�W�tAW���I�I�~q0^.���� �(mi󡆫���7)������>���<�[��jWzؙ��`�%��U�a%sՁV)N��?\.���g�@o�I�rM勃Ua��NN����iW���/S�U�-����	�ɕj��F�c���/T�a����?�j�KB�M@"��S�Z���KGٟu6GN�c�vS��c���AU�2��դ�KM)�U9am��&0��#~w��8_[��U�y�j�)4K�5*\���!:�"<n���̡Q��vj��؂��<�� 
l:���q����c�ꎩ�;���+W��5��S�}E�:��C� ���TDۡqµr�uf�ʰ<��2]��?z2�f�p���8���ܛ����� lـ͸"]�)��7��~�b�m��؈31� ���w&l�e����7��Z�[LS)�4�~�u�V����S��*?e�~�v�^��Fq�ፗ����&�=���}���N�8(w���@���/#_;�l֞U��b0*�tn,hz��Q�[&��@?e��4B��R1���O>���qZ&`�f�%�`e�E�^7Tr�z�g9^E���+宏U9t���n��\�����VD�S21�1��I�?l�D�	����Da�C%.�����k{=Oo]<Rsi�;�-Y�RH{o�����������d�MgO�����D�����l�=�� �|�b��'"�J<�kr4x��n��|%���;
�?�Z�ȏJv�BV�C��ah|��I��e#)� ���J݇s2�'2������>�xݴ���e�ı�89�5���5�h��=�&�ƫh��DȨw�>���L람��M���-^��ތϱ�.�g�Ҹ�Q|+	Ii�'�|1�C���
SN,Ckפxp;�KC�(�����6JԞ��b��2"&$�/�CZ�-��(Ѷ����	��@��K�r�m��������u �����`\"���lX��n�=R)c/�V\|�Ț�dj��3����/��� �W�D�!�g��`��9��H(��h7���,�T�t��c��ˮֱ#j�p� �apػؚ�!��J�dz��_���s�Faҏ7��@Yp{�;�Y"���75U�ӥ���H�Si���n4u�E��.�V�X�$Dr9�*�[��5�o3�(��E��;�c2R�g#�*���}���~Br���I@�W��`��b�L�^���� �c`�?��L�M7Tu�|L��W�B�l4�N�l<���-�:
�f�XD�$Ф��z�q[`lO,*u�߇�1���P&�o8�q)V\녗I6�w�[:�T�U�hG"��i�}��94gݫ$�k�eDƎ�܇���O�4�ڄ���c�/��lq8y�z(����Ώ	?��h�:&����6�^Uxd�?o�,u,��p��X��}B e^��8�7(��Pa-x�E,�n0�ᛛ�+%i���X�Ӗ�.~��W��d&	�G�*?�R厢��Gd���D/W�����0��A7��SϬxޓ�I���z9�Ղ;`.�'�Bɻ��V��g4(t�?\)��O����]_�^�Fc�F�a����&���V��C�lzbp��:�_p��������H����XB�*�).�v���1�*Su��x`�+� yB��ĸs�w��w
4�8�? I=��
��f��V",�q�.\N#�TK�1��l��B�q��X����;���+��[Kt�P�{U���"�?W3� ␐*\޺<�沤j��m�?k�R9!�$`�0ήvjf�1!@�4be�Q	����My�w�G� ;��4�RY��/x����`fO�x�c��T�(O��Y�&���ɖ�p�*�3}����	mc�����{��{tXu%ed:J�0L��@QouV� ���R�<���ۨ�Z��HL�ϵ3ɿ��Hݺ:aE�
�<���6���Υ}�7j�>"���kQ�D2)�J*��4rJ!�/[�MAV!%��_�V0ˡF}��l�������F��Y`��j48�:I��_�+�Lh8��5�]\�����o
�E��!n��ə�w�����U�#�
�9/_W�!�	$'���Q�D�@XX*�g�Ye���{O6�q47�-j|~�`�T|������ٓH.)��O<1� k��I�P(��u������f5�&`�9��]B�aZ?�\��݋P���v��7�KI;R�de�9}�햯3H�6�^�i���zE�pl��!�[��2v蔹3�+#��;���V�9��*Ok�6�j��{%n����Y�X+Ji��G��_\Ϋ�L�>{-��{ȓ��s\*eB��qD�� >u�u��V��MFZl��8�D�̴�(�T�:$�@,^��?�Dz����i�J�q��M�X��=��x�ZI� /�P��%�֑�4j��[ �N �	�t�ǵ��yqWV�4j�.h�%�5մ��
ɰ��_W�I���`�;[�������qx�H��uahиU�e�Y:�/K�%YC�x�B�U�#4�4Z/OHCg�{�tϵ��Y�b^��_��AE��$�/�l�j�!���DF�O7�A_L������j)�a���Xj�]��``p+N!�#[�����!ז@/<��69$�Wc�n@��iEU��F��ѲaGp"�ԃ���>i���������;��J-G#=SEbCɃx��4`O�%P���/-rF=a�����ǂ���>a��;I�r�&���E�1�����D�/*w����Z`�>�^�5��7�m�{G�k�?�	c�}��
� ���л<Tx'ĵU�9�1���_Hj/~k�����/>�9xHr��oc"~���CI��.e��(@�"�����|o�W���5)!M�H}��mr�o�\5_�\11��=[h}�3����`9�c:x:|���"l�#�B��f����7܂�h�ੱ��i�-����P�]��3�|�;!�u\��v9?���g��U��s�ȉRfMH�e�d�Q���j���{����pq�t4І۷�ʊl)�ۧCFpJ�jǷ���˖r5�_���_��R��=�8�x�eUӴ��0��;���S݈P]� 8�z�ma�="�=��|v�T�WMVꢙq���]f��x�w����f�-��%ŧ�T�$Y����dw��1l���d{�|09�⽱c�ܽ�xP�L�7W}�.)̵5�t�����QAW�W�!g��z�+�%Je��H�7\�B��1��Jn�a̓d��BW�͙d�}>� ��4?�_7-T5�.J��"|�pԟ���bK�Q�UF�	��lRYM@ ���7�6�J#j}���=r��AY3�Q^)��Ua��d��h�߀�B/�x�d�l{#)9ŭ�9�4��(�NxJ�/���Ό�ѿw�Qm�u�5bf^����ϕ��6�����2�p K��
3�����P�8R��Nб�l�<��?�4mͮ�/���D_FX ��m$����M��8�����?h:����@9ٲp�ϧ��Qq]Ri�{e��4h.e8$99+�We��A��O;�U��[c�9��nb�y�����K�-(W���v(�|C0�0@�㳩E��&F؈L��M�����Rn��HF���n^&F��=��9�)V�	p�T����Y��*W�/a�z�r���ir�����N�|�{����°�D������ a�7�#�Hqy�5C�ƨ�eϒg��Jy-�m/���t�hU�374�l��W)"�����T߼�z3P: ���Z���?�(UA4{��!	('���1�twɃr��YBG���j��"�zy���Ѻ#�i)�2h!>XR�^��`�,��%B�GIE|��r�?2��EL���-���c�Q4��\=`ǆ��y�?�dʃ�e��J��>����=�0�͋/��5��dp�U�HV�j��D�P���;^�v�BC�`��q�� �3������|Or��>����q���/�iE�w:�����s0o��졏�����TQ �Z[������d��Z�9��(҇<�f-�Wa�m 2��z(�oUhR����A 77<]���HC��%�q�3.�A�T��9lT)�
-�Ӝ����\��|^���nU
&����P�H�ңhy���� ��ǝ�
 ���7X�UGPI7�V�/.S��,A��
�s�Vt�݁w���Zl-�bq���OV@1��L��e�;ue��<I��` $l�"�rv:�T2�%.�l������'	}b!C� ;yE7� ����k�MK�D!pa