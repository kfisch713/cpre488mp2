XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Tg����È�?4�r�XKdJ|-��������<����C��h',y��-/����u���SY�1�Vh��.)=����M.h��Oܐ��<�Nʩ�ϰ����% ���׎:����j9�B_��+�U��_��d(nՙ�(�,����k���i��+���P^�K�_wT� /�.�y�`l���vDK@} ?W���Uj�	�e����y,��aN��
�u�e" ���-�K$]�S��Kz[��J�P�S�Ն��SsBnp$�r���r5oƝ�v���.8�����")��Nd���Zt����TK�#���i*�g�9��A`�=t�x
��x�=��3Y�U;�V�^��ݬ9�+��#M4О����Di�������M���쉰詄���x�)간)���<�Mw�����8�{M���� �.~�D��`p.�I)�>B��r���q%$-��Y�J lp��Z������7,�(����� A����Dml��r[΃���PT�W1t�|�y�qD�lZ��}�48i�)�����ݘ+.�){8�h�iwj�%4-'P:��%~���eh&���kKi�3��IǶd1���!h9D{��س=w�n5����w�Lp�|�� U���Y��������K�%�͓�Vk��853Yd�ʼ��k�I�c�D�^_��2���]�Ⱦ����c1�����]�E�8�묜���h�xH�'��~�@"%�84�w����]B/� ԝ��[���Pc���,�XlxVHYEB    3b09     f80���2Dwa�De�Q���4�\����3�i~EÉ�g>��;T:��*@B�*�G7*�E����&��>��q��`�#����=H����.劇� r�Lߵn8y�0�~�u���1� �'�fo��{;��4���L9"�|L؆�J�Vd����Ɯ
���
*q��
�->-n�䄋��e�u��t�v�݁ג��<K�`Fa�ٗs���n���	"g�ޒ�~ῢ@�3���������,m���)O83�hQ��R����>	q?�������U/ٻ���D��ǩ��ۈ��h
�;���?a?�n��=7T�s�mO+�J�cE����D�k5y�g7�"bNY��B��/ڲ/�l�ڧ�'���ozmQ�kc�[M�H�q���d��~_����bE��?E��vZ�5������-��#�x���	M�ig�[Ux��!�;߼e��e��!�̿ص^�P������z�ʬ�ʗI���4��E�$f� 3�[�!��YƲ��T��@�fw�S��.//����T���VQ�>[ݦ)Q-����FVF����Le�j�2�FoxX��GQ�&q�9��e��i���Jǒ�߻T3A�^��v�
� ��"-�<�Z�z�8��ӣۛrA%Yf<@�Vh��7o�K@����
_G���������d��]������#7�Q(��t��LH�{�b6�)c��|���AJǡ8��z��@�c����|��Z{��������`m6��$��i��f�-!Zi%g 4�%@N�Rd9J�,k1*��~3���y����?�tH{ٺY����t�oނ4��oL6��7��O�iq��-"jv�r|5�����j�gbf<&��X�N�9��@8J~G�+�e
~y��mR.h�&�>��U���s�5|_��	5�_^�s�sB��#fF.���_2�-���(�^�	��ƺj���?�_��&[=��n�)����_��Ruo&\ƯQ�O{#�)3Q��J��@��м�W�[��ީ[c��@�QkOu#"��I���?�>x˯�C�'gJ�j%T�e�U���V��5��Zt�i|�
��l�z�7���I�y*dd�9�O���~ =�l�):-5�014��򐲗-���@�yϴ�)�+`��+�XW�L�@>Wg-��󄬏KF���)	����&q1
E?z�QF�t��G�xh؇�<��,��*��T��x�����M���:Y�"o����9Mj,�
����ߛ���b?�wfc0Pevh-)�+��������d M�+�g�<G'A����Z�>�����H�`Pu+"Ѝ$����GS�H'��T��1���2���,0z�Vƻھ"dٷo)81:QT�
QL*�ʍ!5ǖ�����[����!�:�U��>|A�f�l����N�tR�'�� ֡���ps^�mEpKdbu_���E�$k��W.���8p(�wX��s��DH l_��xD���OM>>���p��cD�����9売�	�����V�+-�@��Z��Z���ߵ��ŋ��w���RZ����:w��
r��k�=�I%앹D͎l4��ݵպ�$񐠕,�ui����q�>��p�J�T�Ar,(>�r)��	�o*��)�e�r�:W�u��t�7Ĳ�~�&cé�i��f!��܌���6Ћj)'� ڑg��WLFŊ���7/A���^'��y�p�IG�G��p�q@��:rxP\�#I�,�
1��jSt	��� "� b���*����=+�gAY���9E���;�������j�Į��۸a�d��j�G���+U��ځ��4�:�n->�������{��h��ߎ��i�������a�^ӿ�_�쏠�nѤ�!�M;2������Z>�j纣Ҭ[�g��Y�	���)�:k}���К��״����7�C����h��#�Qa���B���m�Xp~挙P:��@[F��H$����w(%��,C��էY2������ս�|���	&Ƚ)���7O�����!�S�EyE�q��2�:�.�83C���P5�Te��6%p��DWf�"��Wǘ�=����?�н�oFT?mo=z��Y����`���H�[�\��ijr���z5:$^�a���Q���}Ƥ�]H�!�Tgh�r>��д|���3��_�$.|�η�Ĝ^jX�pw��d����h��`���ē90}p�f b�7�%�.�>/��$�,����<hY�D�x�b�*�:��Ȯ�C����\S:ڶM�������6)i:ێG���"�ꊈGCT���+�w��Q�M>��lc��>���S ��9X��^��ӾX����+(sY��OI��R�	��ou��*��4}��U/:�@V�A�p���h_ޔ�B�<��3 Q�v&"
O/����˔y�'|�p{���4�f�5ϓ��`fd��#�% ���a�=O,JDIl'�C��^vD���NYQ��;*���"x���:�zY�::�8�"�59�qP?��/�C���;�+-or��3:��W>�^�Ɋ�`W܊��̾nX�/��N�{�O2:zˑ�6x�H�ք=�<bZ���v�GX�l��щ���S�Xv�_z��	'�h?�/���&r��C�Ѝ���r��3�Wr`�_vޘ��o-c�N�č�y�c�r������"9w�}
o��l`�[I���)p�L���sւ���֓����卆�6ΩD��D�p�����L�$�_n������7y���k�\T�?�[���4>鲎6K���_��C
`❓8�pX�E����5�ChW�E�lE�C���� c{��Ф@Z=4F'��5���\��R8o ��l��<��۽{�GII��܈0�H���)��O}Q��&6��/�,d�t'�j�6�/���|%���9x�3�G�N�H%<�r��
-ՇU�U�iV�m�^oYB	�4o�]����u���ZiυjJ��<�I������|�dA?/�z34��7-ه����,�;���9�b>�o�o��E����-��8KC�X��s
��^��c[7(B�Iݡ��?��|[,:E�/{�H�Kڦ�b��O�&���#++�=E9\d�y�GO�+4�[�+pR��vN��	�<�G.�����7: �)Db6C�?ErOD�/4�Z�x��g`I��/��:{��|�رym�	�oW��z�`�E�bg8���{m|���VU���wU�)�����9t-]��f����R�X��g1P׊�622�DEg��d h���)J�<�Z�����}�#���;h��.�C�P���l6�f����뇹�`R���z�)��x1�]]�
M(�eoX����c6ĉ���$(��d�C��
�)E/"��[z�&��LE5A�ép6^:�e���L�6��i|�)�'@����C�a�VY4 ���EGԁ�jeZ�Ɏ]Xc2�I�*��R�3���8��$���g���d�T>dWD xB�H#T,�n�CL���ѡQ�a�%>����:@�skU��e��ƋB�� i-��f�E}��#C@�\�Iн�jl�q��j��w,)5l9�J�n�8S����yp������� ���
bT��[�����۹��i/G�jȰ~Xk��f̰,�O!��g�Y��O��-o�N���o2L�X*4�r�9�nr�ajXFN���p�����S�d�Z�C�D�Kv�"&19�vA���I]���Z�F��sU`���	�-۶^q�!����d䡀�{�_q�q{���n|(�n[IS}���&uU�>������#�eP����������,�fw�ۊ*�_Q0�]7D�h�1���B����U�������C�'^�����Iy|0����w���k��}=Eo�F料j}$��oD