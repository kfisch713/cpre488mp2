XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G5�BR|���t�-�x��Hg�X��@ ����
�<�q_��!^f?3 �����=JALg��o]�ᕑ�tӦ�@K$���������t�c��!�#q+$l��R��I't_'�5�V Pwy�8�W��ϡR�c?�O�
D%��۩����ŗ[�;���8[D��R���2�d�� ��������nM��T�5G�^���&I�Te=�ЄM3|��=AT�y�
�]���K�E�GM#��#\����PvK�%�w���%f׾uIp���|��vR��v1�DS��{�R�^��R2�눝�o��O�.H�->6�/S�4�O!iR�+�9�̧��
]�҃���^l�O���c�Q��Y��o�P�9}���ߐ|H�lД����;ڮQɿ������h�o�(&��uĤ?$o��y:<��J��\T�6v:% ����f���~���`R��t�x���Tjg���;,���-j��d��x����,T��&C�u���-U�A��Ѩ��z�*��ѳܧ{5�`b#�^#m�@�reN�AMR��:_���.��f��b}7��)UO� ��E���c����̵����ҝ�kɇs�7lmQ٨�)���YeF>��h��_1�!�?�U����Aхr���[�r5��V�#J/�$Z�*Je,=�u[;�j��3N+�ȉ�,HЂ�J������0��l87��W�$L�k.]��˒0�\{ULL�d�Ґ{RڹXlxVHYEB    3e93    10b0^��cyZ14{�8Jn�S����kD�Y��]x��)���c��x��������*��D���(V[]�:wn�LQ����q�D��pd��p�H��x(��m���_8r⛧[��t�H�I�E���ye�x�!z@T& ����<B����J�4Pg���B��;"W��6c�F\�.Σ�/j�#�X%�q�?����2d)S<9����K�~|!���� ��̦�t�1@�fv��{e9f���j%�?{i�8�st�:e��-Ə2��d�4xHyy��F�=:O	��FSP����Di��j����L��A�����u~M����L��н�����^�`�V��d�����Q��j��0g�m X�]��$�)�C2�+I���j6�!w+�f���3��߷o��a8��\4psA���&��,�<Oc�y�9�-_�i�Ϻ_�=����Vu�@Z���@��P8���?`uX��>�ĭ��}?�έ�U.{w��bI�q/˝�Lv�Z����[Q���,��;�*�����3�a�S&� Z��Q��Ng�҈��-���Es!s�ENTɫU,��J;��vi�v6	ڽ}h�4�ο}�J:pk>O�a~Acitw\�����K���Ջ]��b'U���IQ,gc.7s� �l N��t�$�'����m���);���@���*�Y�8�ە�Zɀk��iBa4B�@"�=�1�8��:;У{�G�i�^�69��/�����3d��U�2,��.��L��_@!2�PG@kw�Gel{]4VX@�Sߍ�ITO��~pn ����EUu/0����)�4F�]���#b�z��N���H��G���?�7��ܿ0'��k��q��E�˻k����>�nP�r�x;u�a�l*nG3�4f���t��x��%��)f:�	c�G���R�,QD%޳څ���vYLc*9�_=�3��.Z�����~�5�Qc$d����N۶�_G���r1�4=��ț0���d�@ڂj��M��W��q�i��;k�AM�a1�g7�Лjp�67����Cܨ �Q2R�a��0Ğ��9R��M:6ݳ�<��D��[�+}�ʣɷ�P�ˊ�[�CZm"9��|�e�V6�}Ļ��|�"�r-�v�I����k�D��zQh�e��hK�]�bѾ�ڞ��I���`S���()�v�de+oҐ��m.����`��D?��-8�}2�?�� ��XF���@Q�◸�L֑(���o;��U����|���s4�e�¸Qn{�'��zȹ� ,���(����L�Oj�&�Tiv6�+��םb*��j������u0�W{1��@�T  ��IC�	�9��J{
�H-������� �4�Ӈ~_�,6HP�{��t`'�j�̌,�#G�1�����%N��7�w�q���"�u���ګ��A�0&aۑ�K�gT#���d/L30nCP9�
��V��ZA����BH���ݓy>�{-��x�2���7Ԭ^�") 4{
_3�F�:�83��ү)�^�u���P{��h�|�.{67x�c�F�[]U]�z����$/&��΀v.A�/-}�(-�5��5fK�����AO�N�"$yk㞨4��!���;�t�-�C"��_8��R����%���9J׬"�3(q+�
�� �k�hk�����K� ��ƿa����	�	��E�vƣ�=c'	k��Tb��)��<9��|�������߇S5ie�z9L�����ުx{�ZՒG��|�� @��Q�!�(������:M���DTL�W$z�,B�����D�^m���GeΑ�[}01�v�jX��FX�IV�K��_!kf��6�����fT�Rȼ��Y��Cd�߶&�J#�Ij���L�׫���8R�w���@#��A<�O�lM1�n�/a?�"��8I!u
����3�t���}N����>�@������T�B��)<��Ê}���W�+)
�赳
')�W�����u&<������'"�r�E�c��Zx���}1}JL�sd��G&�=ys5��۴��$�6�q�p_�s�^�?�M���D����\���^N��z.7����r��.H;=2(����T�d�̫Vĵ��8m������ Ӂ1�:o�q\�`t@P���x�S��L]����5��!R2%�PFn��TOJ5q�f>q�/�jx{��"Q[vx�t�=�M�� �[�j1�I�K�|��T�Ȓ�W
H��1wdn�a2]��"�غ8cUj�2�&'Jf��S>Wb�`/P��q#Toṇ�z7��t+oҁ)Z��5���R�S�껕�NB�uR�	C��L0������FR�	�Cf}���\��BN[�ok��x9�HXp7� �'�#H�2������&*-�=M�uI���U0)��s�m*Yht�1����{|{���S͖A� ���Q��9��G���Z�v���=��oH�Ql��S��P:x_ ��$^�b�H�[����f��MC�1=l���V���̔w2f��ßS�7F��
OF�4&��/�D�M��֯c=k �R@v!�\i��x!Esg��:�wA�XUO�l�x���#����e`�SD\؅�b�_��EД�i�Ā\j���%��? ��\��&�ֵ�^�@����U�µ�@6Յ�g0�1��	��]�EZ˕M|�m]��T@n��ׁGЏ��q
r��A�*�&MsR-a�laq�$��D�����V5in�W
3�nN���y����U@�rJw>+��X������;��e1:�&iO�>���Nl����OY�k��O@���Q����']��]�,�k��K��`2e'��V
M����s�|F�"^��%Ӹ��)Q�Op�)�"i��HQ�~��d>�"��1DT�ȴ�D���X��4���x:S��$6 n����he3����T�q�c�C��]��%@i��`� ��M;�WWR��V�t� ���-j.����b��αp��a��1xfR�����hG�*gt�8��Ǿ+x�m`�U�cvosԝ��XN��vI��m��?(-�l謖ߖ��s���(�܂�"���㐀���Hl��0E��]>R�&�@��ĝ�����$k\�4\��z[b��iG4��}�)�U���(�Bv��/��?57�9Y��%;���h4����0�5���ȜZ�Ya�<�/� 1��6B��qt��~-�j���R^�Ū���@�zfD
�ɰ�[�U����L�o@����Nx�.Jͷ��D8ʓ��H�?����i�=���s�]�*�o��p^-���T�7z���t۾�e|�1�yU�F�>�i�@�P;
NuR������!?Nݛ@Vg	��oL����̈ӏ�d��T�]P��`��ԕ�=�oiBQ��7gl+�]�DYn��\�9ݶy�����c��k^���b��I.�4/S��//�H����:�w� ��K휍a����k����B��]-�-�R�G�@!U<���G�j�3L�l�3���-$�L�o/q�k%���#�/x11��Wi��� -ȷ��4Q�`!�]�dؚ��׮Vټ�i۱�'����,t���O&ݜj�"�����I0]{�.�e2'�%a{#��(GX͉�����K_Va))�qF�Ql�%Ӯ����65B�E��	��F�����ڃ�{��[�T� x�a��	�B���D�^�Z<#nF����M%�����֗��g{>�n���J-:�`ŝG���Dᰑ���#S\�����}��%��=*B�����H=�0�$���|D�S3u)l�a�R����n%"��ܙ&�Jm�Uw��b���b�@@3L�ӕ�]Dw��}����?O �������[���3�l� n��9=!�.���+�@}�� �?�!�9H��i|H�T��zh��y	�y��YxtI���{�=1����β������j~��"�×���\�`.�S�MF⬓-!)�Y�n��;Hg��<���&��#�1KP���d�$#a�@�WU��L�t�U��m4�Œ::�Œ�U8Q�`����}��(^0Y, y�6t��K����8�'b�L�ݧX?�ȡ�x�����Uݏ,��Gz@L�����q�4a�z��}�,:����~�N��'ܯ��{=&���w�����P�����͡~�'�]R���F�3�!�)6�m�Y#�P��7�S�%�����iMs�o1�t��p��W�4�[�-+��-���P*o