XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��aq�_���c�~8��ķ��pf�nQ�������Q��p����{���1��]��D�A\,t�}�:̊+t)���B���<¸Ye�Y���m�]:a)���?@ðO���^dn;,S�Il�I��z�m$��=t������&R���k�z�o!E�Bis/ �v?�ŰQ\oL<J9�Ӭ<�q�ҚJ5���*<UF^����D*�ك\��#	���������تc�5O�=PٴE�!v^K�h���
E��&��n�=��k�����[~�1o�f�5n,�ȵ�������k���žj�ZZ��jC?��@���s�x��
%^4)��׳�k�$��ʈZ��>7*W�ׇ�Ř�a�%�+=�f(P�E�R���D�&��|G~��D	>#Z��N�-�P��.c�gB ����R[|�^D�{�mR� "�s��|b���lw.�M�ޚ���"�J��C��N֟7_Mu(K!�C��C���USeFC�NP,!g�!Dԫ��Kʨ��=L�����ڈ�g��.E)��P���'��}2�00(C�>����u.�i.HL�T|v�?/.��k ��v4�/E2m�Ε�� D����P	9��ȹ��-��h$w�n���	!!v�E���$2mJ⥒<��/��\� *���uP�y�u�oʈO��j60�F��I���yXG��O�!b�&��H�Kb�r��G�%+��z�y`�Z��J#���B�⤑T��<Ye.�;�U�IM0�����8UŚ0NXlxVHYEB    374e     ea0��$��Pq��F�"�V��U��-���"ƴ��{S��8���D���/���N�Clt���jd�P��ܯq6�{-ϊsS8 �/�e��@^�3tl���BƗ"=0�h�Ƨ��A+8@Z��}�'I���eaP�~%ʲŸ旄�d���c��#�~�E D��`y�Vy��L�\W����S;7,�L�hp�,i#j8^��v(�E�\���B� x�Ģ�Ǥ���tB���	��|���<`I!���9#�w��*#y'�c��!��vGǌ+s$�^��
�-�1��DG��M�i��E)�����k��SY��[�������E;=F����x���������u��?@a�zb�T��s �7�yh�o%0+���\'�?^����Y���15��E�/%0**�?`m��N�0�S���Y���p�������]mL3��N8�C��~$R�Gp3�cc�'/#}�r�X�T=��z[;�XT��;Ƒ3�s|�T��^KtQ7d��������d�0�e���2�n���ݏ�������[�4vx잁,%�ce�S�W�ܸU���>,bt�����*� |5/�Yc�5��=�F_ryӕ�}��t���,j�s�p������]B�9"�f����_Ŋ�v|+�1�0z'G �����y$�N��Ť`
��]�J$�E����U�U2TM��ws}��Fa�'�D�:���ŗ�D�jo�R�xS� Tɔ�,%.�)2'��`�h�j#,Ξ�0B�u]�Q����7��:y1�c tjO��	�-��K�|�C�L�������mZ?�E4���~K�A��|C!1���ŊH��^x�nġ����Ǽ>���G0q���e� ����c���k�m��,�(%3q��z{Za�Y���\�T�}�X@�����_���NT��^PڐY5'1~�K����jBnIʙ8/Sv+�h�K�c�����J�L��x�DcFYY�]�H�qU�������j|-(O�kh�0�^�6�}�u;=$đ�Q��	N��n������9��R}o!�t�����;5���+tf��4�߻���Q@��ef��;r>lu:C�jdn��E�������`%]���H^�Z���]�x�wi �r��'���T�i񥾳����b��u*�� cBo��AZ)�ss�:J��1�pU�����a-*�eL;��q���b�������C��[	��*���Ui
c��zf��+��z'�@�eP�rMn�#kK��"Rd ��k��I��PkC	t��I�� ]�>k)��$\,`���#;I`��~i3���*��l�X�透']^�:C�Zp����L�K��^��ٳ[�t�Q���cwVb@���B�a6P�e#+�#OY)�=JP\*+�X��` �]b�����������|J$:��w��:��q���{�N�/��������]u^ﲩy�=�9������*��|�I�>?"� ar�����0�||Q��ر�/��[m��,;��q�3��m�?o s�#��(GV]v�Q/j���8�u�*< ��O�����[���0l�VN�/+b�������d�7hKkv��И�[	e0w�y��.%K�D�E��/_�����]�����ԦR1���̢p��G��d�/.ň\lPכ��ގ�j\3��|"Ee�-�"'U���#a�&	H*�����&�@��������݌��*�IRP��.jE�ŐiB���5�� o:@��#�A*H�aA��	S��IӍ�~w��w��/���L�7Z�<���v��d^l	�BAJ�2���B�O�?�7zt�����'ƪ�/�Z�D����Y?�W ���[�d:���yO��b�(d�����l���G�c�9]T�s>����7���7{��l�O������0.PЗ�x�S}/l	���y!(~��:� �}\�޷�=����N��>g�SR4�DE�k�zNmF��mՙ{���N��ְ���G������d,�i|l�P�؁Dտx���a�T�9����P�_��k����.�U$�|e��-��]TB[��2�����7r��mnZrzh����Ӽn|�N�C���,�V����˯�	�<P�6��ui4\��z�PːƗ�Aa����u	�E����ȭ���@��c��SЎ��!?)��X��W
f��-M�в�� ��A��I�D\����ᰖ�Ti���/!���8}�6Q�qxJ�ʑZ�7d�#}�_��xFm�BD�"$9�F ������,���.鬌�Z��I���~�g�_�w'�������u�BÙ/��B�
_"4Eb��p�ܩY[�p�> $_S,�9�:�������Ùh˿����-[�l�@{���a�u��g��4���2ԕ��`p둽�2��V�R���dT	E����p�:�p��!(���ur7��~�+�k$O�!�Cݛ�!m��K3�_Ps��t��mt��fw;{���:�# 1�r#v��/Gw=��o����3�M����;}��n8;Ә���~6w]ު%���f/�S`�oF�NCa������O�`�u���hy2�K�&u�XDp�t�X@�Cz�֠��\Z�c�!�d�j	�dw�����W4pAiE�w���WP�æ矤w��vd��9���6�RL
��(]-� �) kJҏ��o=#"��>�9���'UR/��O؜��Z|(�Y�tΐ_�@����C~��Hl�bE-u����g��6���	���[��kr��T,�軹*Z0y�n�Y��.MK	�iz8I��ڮ|5'xl{�U�1!>�;+B��e�P��#+]N��ָ�E�ܓH�uˠ�xE���B;�a���A�ks�	J�Մ�䡖 5?���t�:9$�!'�ӿ�����Y�f����Y.z*�eU�XS7�O�gC�Ž�oZ�=
��4k��n�-n	6i�_5�㚤^�Z`��T�!�kh*źo�R�hC��.�?"~�t���,����1�8�N��}=y~����2�Ǫ�I�^��%�B�,�����{+����F�`�z�'���̙#��`���L,:�Z���ͧ!���M��}���o��W!�`���:����ֶ�sM!v�g?��Gc�j>cq�C(]�q�Dړ�|W�5Z��Y���
��Q��J4Y�1?j{Gˑc��I��9׃�Y������K�}T�J�p~��inD�ͺ����Z����'> �?��iF{�v�ʪ������\�H�<��E���ӕaT3�)����k��˦�S( ���3��xs@��Ƨ�����:6�	�g�6�ξ��cV[ȏ��|Bo�� xn���&����'4hY��0Cǖw�/A`~s'8r����B+[SxT�(�Sf��8�-��Ĉ"��l�d�鱰L�$	̫��b�r\b"������ɠ��Dq+�U+���3!3�����q�{?shU'v?�F*ڴV�5�#��,��R��W�gݱ��cq#xU������j�{����T�#l�F�\�!:�WY܃��<G�!��I�8����>�"�!����M�[��G�f�gĊw�bmE��� � ��L�!n�򘅯<)VS�qC��Q��e��I5c�aލ(�0P��r^0�j-�6z��x��j���-I��]*�7�\%P@����i� �p`v�