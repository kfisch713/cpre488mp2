XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��fK&#�s��$P�(a�T<��љ|��}�Ni*��9L��\�!Ov�?4�⹩&S���86M�T�,W�9�P�Uq�?�!���k/ A�I�^��J?{j؎>��~��4鶼$�G
L��VP4A��}�H�V���x�OQ���V���oҬ�����Nh_>e#vH4��T��0�Q��u���	�iwA]~� b	����&�� ��
������Q�f�ڊs�7���^5U9 �?�I��^���(W�zI�"��Bf� C�"�.CX���	�y�5D���;�� l������\�Z�'c������槢���)oJU�Z����H ���V�c�>f��f?��yZOW�im����(5ޙe��d�\VX���.Ņ��ï�r���f"�*�6��	ad}��.�̟]v�+�;���t�bȃٓ��(�4����_�!�q{߾����o^����jg;>!X��t�<��P�a�yw"�\�=w	7EG���W������L���C	�ۜb��@^O�9��w�X �ڔť�3Z{�P��d#�,[��K��m�l%r��ً�S��9��8��vu�L�����}V��~|�C����w�$$:��.cK���C6�t}��y��a���M:{��5ۢ�/��h,��.qI霒މ�u�DE'�%�I�3�4�ݕ)�@(���#���g?��T�9
*�u�l�v�0.#^y�G*��g�)�^AՋjNGY<x04 �wEUz���@"�/XlxVHYEB    290e     af0nw�H1*;/Qw0$�å����������Uh�u��>\��i�ֈ���c@ ���ѷ���o�K*�n������%OD:���s5��G�_>�j���z�#���U���f��K��_��v2��#S[q;N��0n�Ʒ�b6'��޹��'3����{��!:0�<�	O_~��+�t��>ν�m썤��A&�D�-���Ɛi�����e�
�E���J%ѿ����~�����[*�%IG����5k�B����5Q{|\	tV�qĚ�z����M":;g��Z*MД���;�X5�4�[�16 C�kƘ{(	S��jz�w��J���Yu�\���'�Eq��RE�hy�r��ݕ[�Y�6������Sh�'�� �ˋg�%}��W����çˀ:R�U�����?~>�wwEm�U�h�:0���=�b��<I��TpC��*�x�a���������U|0�~�@��qϜ<����ۢu��2�@�ʰ�Ӯ���K��ZS�o�'�'��&�ؗ'��/� t��#0��)8�MxrzRL8V F2��'ƿ6>h�3�B}�X7�0�_��:��3-.�Ud��q@�R�Y�𛢔߂>��M���\Ue<�����͖[�@2�"�g����l���5(����Z���gz�>�I�k+���|���IV/�&��߿~N���iv���R�KT�A�X�����<!Ŵ�y���q�?
��z�rb��G�f�Ro��r�/߾N��!œ�/���.��^�\)�"�Qj�Y&�-g�MI#G�c��r�;ڴ_���	Hy���������*r6%VN��a��!��XZK1����S�p���&Y"�\)1^��9}��׮�5��ɽߖk�lm�`F�y���Z������f�(� _u�D;�ʋ4/��.�5M�^p�����@P�K�Ir� ��^��x�m�7�9��[�� ���~N�DK���|�w�'�<��h��5��F����>�����v�J��p�EH)�a!��0�C�s��k�L��rݲ7����@#�劻`�zl��m?_��)i6g1ȳ�n�~��4���A� I�3V�M���G��TZ�4���whc��l*���j9��.e߆@L���?��� �������¹�zx�~��&D�=�{���i/Q҆c�Nl2�O@����i�#�������su3��Q�/z"���|��� �� 3ݬ2�"ߖm[&����Ṳ�9b"���<��O1���"���-C�E��S�P��=���üIM0��h�m^q���+�-#�
�����%�G������3R
���k�Θ�ͅD�׿(%h�#d9ǳ��v�� �	(�������@��ǭ9 ]Kx��}��t"�;���8�N��~���+�_zz'�c�п����f%a�K�C��P�tf8�s�ˬBƴ�N�x�a���d�Y��C�UB&�YG�����م>��.GNa�^���c��`�!�)�}4e�.�a66|A�+�@��~������%��Sے(^�⸚�t�����%F��1Z��ΡS���Qt�^Z�U6�?U�##qӤS���
M��٨#�Q�tW�ِQoב�+���t���_�P�%?�l�T��@�P��x/3���w|����nW���U+�`4�j&��[�A/��l%D�!Ar}{�Ҏ,�y*T�v3]���{����=�}�Q������E��r�';�P_���U�A#8a��C�^x'�_��A�I��#��ԧ���&�}	�qs�}�/^�tJ���)�B�D�I#�P�m��Oce�5�L�D���x��1�o��tҮ��Ӟת0���>VDǧF�7�@�� ���C����K:n��<�9��,4a��3Y5��qjx(��^Hp�,c�vl<�!��5U!��fo�#�%�d������+�4R:M��@9q$i��i�H�F#�.�kJ
��j$["�0g-�T
)9�ϧ�tC�z$C���\���k f�f��Ǣ�lX"��C�q��.9�H?<!�-��x�,A��f����.Y���Esw�j;��:�"�J���;o� ��������S��:�톷ǁ��J����Sm$N��?K�kP�f-rg�s�l��j�뉲�Jts
`W4 3zF����C�����ۃ&e�qo?�*?�ֺ�YQM+<�)#���L��\��Z�S��c��7@�"�B��fhTu�>{c��z���j
�5B%���n2ʗǙ�a�DY��:}&�s.�=������n����'5��V��`�~���ޒ.�m�7>��Fx���BV�Zj�IVZ�勂���܄�{dk���J+c�~�7f�%��Vv����i��pX�g0�J�k��}-�{��ū���*Ԇ���䏏�W	�c�GJ�FN���HPhX�*���?��i] �
��;�����o%M�������,e��_��=�š�q�	�R���F�+6"ֱNdգ�@�F���Ii�mMo��;]$��BVLW��u��M�y��icH�&E(�l�5X����G�&Lw��{L�1-� �PT16zd��3o��!Hw��ɛ�r�)�f]dS�Q���pn�Gje�&��)gF�� ���(�	���5�|د�饫��P�G�k%����C; ��8'*�ؗ4��c�d9x$���5�>��&���:-��7)�:�o���+�+����*w�^�
'���8��N������{Uۙˤ�z�z+�n�@t��oږg}tsn����Ȼ�̊o