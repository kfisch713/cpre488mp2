XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n��1~����/��rM�
"��	�_i�T�l�B��tA����L�y��e~U����6���y�k8�����u(w��aH�9��{��}��{�*u�ͣ�^c�z�{ď뿬e\/�4Q̨&��w;�Lnb�fwĬ-���j��z��ħ�E��tc+��c��W@t�C�t��1:�D�#�M��(!^r��U�/�O|*7~,��D�����T[��?�?�Qtqv��ɉ��S|�)K�9�n��>� $!��}6!���v�/t����-/����Q�}$ ߾6�2�"����J��9�h�W6�!�Fݐ���R%:�9�W1Cn.�Gxb��D!?�ӻ�6[���@���n J?�s�\b��f)Z
� ��>Lu��A�-�D�(��Q2��J~�Q���9�Nt�L��Q^q�-��"��lF�K'���;��ek
#���[׵m�d�F�Fd�?T����S	b�t��71����xP؎�!��\I����M�	�i|U�vYt^�B�(��Ȳ���MN�%���+���0|@��;��"M��=8����������yhz�]�jճ6f����yAd�I���$��J!\� ��x�7-���G�b�"���5�����,`x�7sϺ�0����D:>u�a&0>�d8����y�!7�P${�i��O�jf�XJ�n�݂ο֏�SA]�-��^��jf)��e�����T�W�W�{���|�E��q�n�D )��{y�5�<�Og[ᠵ�e�Ԙ��XlxVHYEB    1a2e     8b0&�������U��?&pt�8���zIT"vbIE��XkӲ�Z�@���fg�Q����[bfiNܾ�k���Q퉵��SҩV%�7g���ԚrqX��8&u�H9�N�����e�`���8����Q���GV���{�m��S�_�MB3{v�;�du��1�^��o���ωJ�*�%�b��+�b;�P�u��~V=�ǦoD+��/t<F�uq�<�(�S��zruk8�~)n[�}\���ΡU%�ޱ[���M����L����uI��Fdq˓��cz��{�{�IGOh<�}1#=�ˑ��B�O7��]���|xp��L������Xwf�	���B��dK{�=6�$Q`[c\�z:��$NX�>��:�,s�9����bŴ\W��b���ؙU>���EW�g�3wC�����z����+�dZ5��M_����צ{F��G��~7�7(�������7�t��r>(�
<��gng�^n����C�˒�XM��wA��y��7�/����+ZP�������5f#D[�ٹa=to~�Q��5�;��~]Ɣ�2��-����\� !�LR���4o�M}v��I��. �f��.�I/�r
DXK�M>F�l��Ɣ������ބ}㤐U��H��4�D�!����<ȍ�,`5c��J� zL#�����P+�m��� ��_�%�׿��?l��z�S�߁S��I ���ނK������3�i$���qDJ��:y�=eK��ԛN@�E������u�g�_Gj�k̠B��K©���4��.��ޔ�`��hx�2;� ^�(�P�����[�1z����)�Y٠�[	�R��5�cE���O^��G���bW��U@��\�j���#���G)�m0�S��~O�{�"IQ (�.���pԣ8$��?����lXk�i�QL/�~��3Y��z����ܲx#���̗bg�|_��Swd@��!�s,'���󧋶�ThyZ,�sϳ�����q�87���GA&���J���H\ﶣ��"���'�妪��<���W���������]((�>�j�ߦ=�w�l�`t��0'�����`�cdP���O蓼�L�E�-^�)�����a������P�2��,fRɓ��y�Ugn��j�[ThZ��D/ΙB/���TU�o�>4�_�v���Z��f����A4X�#����X$�(���X�U~M���� Up���)>j������=�<�δ(���
��2��0�7D�,���}�T��lt�_EԥXx�>�P]�Xbօ��&-��T��oS[y�"hYe8�t��OqY�Kp�D�W�g�pȲ�A�[��ָ�{�&a=�b@�y�}%`]˹%������z�+?�����^
�N��}"�CjO ���tH�� cJ#���`N��C3��J�D�ur��m���<ح^m�bJ��,.��8�z��@�ڝ�"X�}i�EN�~��+�G���s��~%f��
�q�y��S���dOyu�}���L����O&������{�"jM�c\�m�xV_#��[��T�k撗I٬��q{�Y�����wi���vky,�2mA>E?ݮm9�O�����;.5ߤa���WK��Pk���Y� �!�a�ۣA�m��7��L4ʜ��?�|��Py��,�P&ҏ*���C;���R5�Ɛ)u
�t�������E�τ��쳀ރ��t7�gӘ��	M���#+f2��Jٵ�|��K��$�PШ�~qL��g�S�f�d���ĵ���5P��ۡL_vxժ���1D�0���myKǳ@�P�Po*���m���a�D�A�Æ��>#�Ӂ��!,����Ͳdm���,�쿅#�� �t�`A��B�-��1�R:Y+�P&Qe�����*��O���W�W��1��X�P��	�,@3J�n.���?�e]�����
̱�;vF8�IҐ��6�č�&n��Mߊ����=gC*6�&�o��6:��tJ=j����,_/����y:s|c�M1g
����,�M X�.Y%�4�d�	=��#{LQF�̺l�S�����t�s�Ӧ�u��7@�8�/�8f�G���+	W��H�$yF��mE��,�6�O�%�˾�����Vj��!�	�\�i�H���dh�z���h��m�X�w��E���*�P��o��`